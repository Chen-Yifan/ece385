---------------------------------------------------------------------------
--      MassiveSprites.vhd                                               --
--      Matthew Grawe & Larry Resnik                                     --
--      Spring 2014 ECE 385 Final Project                                --
---------------------------------------------------------------------------
-- MassiveSprites stores all massive images.
-- Namely, it stores the title screen and pause screen.

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

entity MassiveSprites is
Port (  Clk : in std_logic;
        -- The row of either image to access. 8 bits because 2^9 = 512 to reach row 320.
        -- Well, one bit less would've been fine actually.
        -- Addr selects from both Title and Pause screens simultaneously.
        Addr : in std_logic_vector(7 downto 0);
        -- The color bits of one row of the images. 320 because the images are 160x144
        -- in dimension with 2 bits per pixel. (320 = 2 * 160)
        TitleHorizontalColors : out std_logic_vector(319 downto 0);
        PauseHorizontalColors : out std_logic_vector(319 downto 0));
end MassiveSprites;

architecture Behavioral of MassiveSprites is

constant IMAGE_HEIGHT : integer := 144;
-- Number of bits needed to represent a pixel color.
constant PIXEL_SIZE : integer := 2;
constant IMAGE_WIDTH : integer := 160;
-- Number of bits needed to represent a row of pixel colors.
-- It equals the size of a pixel color times the number of pixels in a row.
constant ROW_PIXELS : integer := PIXEL_SIZE * IMAGE_WIDTH;
type rom_type is array(0 to IMAGE_HEIGHT-1) of std_logic_vector(ROW_PIXELS-1 downto 0);

constant TITLE_SCREEN : rom_type := (
x"aaaaaaaaaaaabfffffffffffffffeaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa",
x"aaaaaaaaaaaabffffffffffffffffaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa",
x"aaaaaaaaaaabfffffffffffffffffeaabffaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa",
x"aaaaaaaaaaaffffffffffffffffffeabffffaaaaaaaaaaaaaaaaaaabffeaaaaaaaaaaaaaaaaaaaaa",
x"aaaaaaaaaabfffffffffffffffffffafffffeaaaaaaaaaaaaaaaaabffffeaaaaaaaaaaaaaaaaaaaa",
x"aaaaaaaaaabfffffffffffffffffffbffffffaaaaaaaaaaaaaaaaaffffffeaaaaaaaaaaaaaaaaaaa",
x"aaaaabffaafffffffffffffffffffffffffffaaaaaaaaaaaaaaaabfffffffaaaaaaaaaaaaaaaaaaa",
x"aaaabffffaffffffffffffffffffffffffffffffaaaaaaaaaaaaaffffffffeaaaaaaaaaaaaaaaaaa",
x"aaaafffffffffffffffffffffffffffffffffffffeaaaaaaaaaabffffffffeaaaaaaaaaaaaaaaaaa",
x"aaabffffffffffffffffffffffffffffffffffffffeaaaaaaaaabfffffffffaaaaaaaaaaaaaaaaaa",
x"aaaffffffffffffffffffffffffffffffffffffffffaaabffeaaffffffffffffaaaaaaaaaaaaaaaa",
x"aaaf0000000000000f000000fffffffffffffffffffeabffffeaffffffffffffeaaaaaaaaaaaaaaa",
x"aabf1505555055554c554155000000ffffffffffffffaffffffaffffffeffffffaaaaaaaaaaaaaaa",
x"eabf1505555055554c55415550555500f00fffffffffbffffffefffffffffffffaaaaaaaaaaaaaaa",
x"febc9919998199998c99815545555555055003ffffffffffffffffffffeffffffeaaaaaaaaaaaaaa",
x"fffc642666426666426646662666655545555403f000ffffffffffffffeffffffeaaaaaaaaaaaaaa",
x"fffca8aaaa8a9999819989991999999919555554055503f003fffffffeeeffffffaaffffaaaaaaaa",
x"fff2aaaaaa0aaaaa82aa46646666266626666554555554015403ffffffabffffffaffffffaaaaaaa",
x"fff2aaaaaa0aaaaa82aaaaa899981998999999919955554555500fffff8abaffffbffffffeaaaaaa",
x"fff2aaaaa82aaaaa0aaaaaa8aaa8666426666662666655455550503fff3fffffffffffffffaaaaaa",
x"fff19999982aa2aa0aaaaaaa2aaaaa98001999899989991995515540ff3fbfffffffffffffeaaaaa",
x"ffc66662646642aa0aaaaaaa2aaaaaa26002664666066626664155553c03ffffffffffffffeaaaaa",
x"ffc99989909901990aaaaaaa0aaaaaa2aa99998999099899998995553c03fffffffffffffffaaaaa",
x"ffc55505626642662666aaa810aaaa8aaaaaa64666666466664666548000fffffffffffffffaaaaa",
x"ff15551551599999199999980aaaaa8aaaaaaa02a999989999199990000003fffffffffffffffaaa",
x"ff15541541555666264664606666aa2aaaaaa0a82aa66266662666000000003fffffffffffffffaa",
x"ff15505545550155198998899999990aaaaa8aaaaaaaa199999998000000000fffffffffffffffea",
x"ff0000554554015455066026666664000aaa2aaaaaaa8aa66666600000000003fffffffffffffffa",
x"ff000000000001545515509999999898009a2aaaaaaa8aaa9999800111000000fffffffffffffffe",
x"ff00000000000000551541556426626666646aaaaaaa8aaaaa660006644000003ffc0003fffffffe",
x"ffffffc0000000000015415540599199999899aa8aaa2aaaaaa90019991000003fc1555403ffffff",
x"ffffffffffff00000000001500554556666466660aaa2aaaaaa80046a54400000f255555543fffff",
x"f0300003ffffffff00000000005545555598999909a8aaaaaaa80019991000000c9995555543ffff",
x"f2022aa3ffffffffffff00000c0005555554666666646aaaaaa80046644400000266665555543fff",
x"f28a0203ffffffffffffffc03c00000155545559999199aaaaa000115110000001999999555543ff",
x"f222323fffffffffffffffffff0000000055155566626666aaa000444444000006666666655550ff",
x"f202323ffffffffffffffffffffff00000000555559199199aa000111110000009999999995550ff",
x"f030303f0000ffffffc0003ffffffffc0000001555466626666000044440000006666640666540ff",
x"ffffffc05554fffffc1555403fffffffff00000055455899919000011100000009999901999943ff",
x"fffffc1555553fffc155555543fffffffffff00000055466626000000000000006666602666603ff",
x"ffffc15555553fff15555555543fffffffffffc00000505989900000000000000a99998999990fff",
x"ffff155555554ffc55555555554fffffffffffff00000055466000000000000002aa666666640fff",
x"fffc555555554ff1555555555553ffffffffffffff000055059800000000000aa80aa99999983fff",
x"fffc6666666663f2666666666664fffffffffffffff0000505540000000000aaaaa2aa6666603fff",
x"fff19999919993c99999999999993fffffffffffffffc00005540000000002aaaaaaaaa99990ffff",
x"fff26666426664c66666666666664fffffffffffffffff000050000000000aaaaaaaaaaaa640ffff",
x"fff199998099980999999999999993fffffffffffffffff00000c00000002aaaaaaaaaaaaa03ffff",
x"fff266664066660666666666666664ffffffffffffffffffc000f00000002aaaaaaaaaaaaa0fffff",
x"fff2aaaaa02aaa02aaaaaaaaaaaaa8fffffffffffffffffffc03fc00000019aaaaaaaaaaa80fffff",
x"fff0aaaaaaaaaa82aaaaa80aaaaaaa3fffffffffffffffffffffff0000006666aaaaaaaaa83fffff",
x"fff0aaaaaaaaaa80aaaaa000aaaaaa3ffffffffffffffffffffffff000009999aaaaaaaaa03fffff",
x"fff02aaaaaaaaaa0aaaaa0002aaaaa8fffffffffffffffffffffffffc00066666680aaaaa0ffffff",
x"fffc0aaaaaaaaaa02aaaa8000aaaaa8ffffffffffffffffffffffffffffc99999902aaaa80ffffff",
x"fffc00aaaaaaaaa80000000002aaaaa3fffffffffffffffffffffffffffc66666602aaaa83ffffff",
x"ffff00002aaaaaa80000000000aaaaa3fffffffffffffffffffffffffffc199999899aaa03ffffff",
x"ffffc026666666660666666660666664fffffffffffffffffffffffffffc2666666666a80fffffff",
x"fffff199999999990999999990199998ffffffffffffffffffffffffffff0599999999983fffffff",
x"ffffc666666426664266666664266664ffffffffffffffffffffffffffff0556666666603fffffff",
x"ffff1999999019998199999998099998ffffffffffffffffffffffffffffc15599999990ffffffff",
x"ffff2666666006666066666666066664ffffffffffffffffffffffffffffc05556666640ffffffff",
x"ffff1999999009999099999999099998fffffffffffffffffffffffffffff01555999983ffffffff",
x"ffff1555555401555415555400055554fffffffffffffffffffffffffffffc0155566603ffffffff",
x"ffff1555555501555415555500155554ffffffffffffffffffffffffffffff001555990fffffffff",
x"ffff1555555555555505555555555550fffffffffffffffffffffffffffffff00155540fffffffff",
x"ffff0555555555555505555555555550ffffffffffffffffffffffffffffffff0015503fffffffff",
x"ffff0555555555555541555555555540fffffffffffffffffffffffffffffffff001503fffff57ff",
x"ffff0155555555555541555155555500ffffffffffffffffffffffffffffffffff0000fffff555ff",
x"ffff0015555555555550555415555000fffffffffffffffffffffffffffffffffff000ffffd555ff",
x"ffff0000555555555550555501550003ffffffffffffffffffffffffffffffffffff03ffffd5557f",
x"ffffc000000000000000000000000003ffffffffffffffffffffffffffffffffffffffffff55557f",
x"ffffc00000000000000000000000000fffffffffffffffffffffffffffffffffffffffffff55555f",
x"fffff00000000000000000000000003ffffffffffffffffffffffffffffffffffffffffffd55555f",
x"fffffc000000000000000000000000fffffffffffffffffffffffffffffffffffffffffffd555557",
x"ffffffc0000000000000000000000ffffffffffffffffffffffffffffffffffffffffffff5555557",
x"fffffffc02900000000000000000fffffffffffffffffffffffffffffffffffffffffffff5555557",
x"ffffffffcaa9000ffffffffffffffffffffffffffffffffffffffffffffffffffffffffff5401557",
x"ffffffffca905553ffffffffffffffffffffffffffffffffffffffffffffffffffffffffd52a8557",
x"ffffffff2aaaaa94ffffffffffffffffffffffffffffffffffffffffffffffffffffffffd4aaa155",
x"ffffffff2aaaaaa53ffffffffffffffffffffffffffffffffffffffffffffffffc00000014aaa155",
x"fc003ffc06aaaaa53fffffffffffffffffffffffffffffffffffffffffffffffc2aaaaaa80aa9155",
x"f2aa8000016aaaa53fffffffffffffffffffffffffffffffffffffffffffffff2aaaaaaaa80a5155",
x"f1502aaa0015aa9417ffffffffffffffffff57ffffffffffffffffffffff57ff2aaaaaaaaa215155",
x"fc5542aa8001555455fffffffffffffffff555ffffffffffdffffffffff555fca8000000aa814555",
x"ff01542a9000000055ffffffff5fffffffd555ffffffff5f5fffffffffd555fc815555402aa01555",
x"fd581282a4000000557c00000000000000000000000000000000000000001572802aa8004aa15555",
x"f5568aa8294000001572aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa8572200a800952a85555",
x"f5568a800aa40000154a0000000000000000000000000000000000000000a152282aa82a52a85555",
x"f5568a01506a00000528ffffffffffffffffffffffffffffffffffffffff2852282aa82a52a85555",
x"d5558840251554005023ffffffffffffffffffffffffffffffffffffffffc852282aa82a52a85555",
x"d55588680a4155555503ffffffffffffffffffffffffffffffffffffffffc852282aa82a52a85555",
x"d55528682a9001555554ffffffffffffffffffffffffffffffffffffffffc852282aa82a52a85555",
x"555528682aa054001554ffffffffffffffffffffffffffffffffffffffffc852282aa82a52a85555",
x"555528a82aa050080003ffffffffffffffffffffffffffffffffffffffffc852282aa82a52a85555",
x"555528a82a8005480523ffffffffffffffffffffffffffffffffffffffffc852282aa82a52a85555",
x"555528a80020a9484123ffffffffffffffffffffffffffffffffffffffffc852286aa86a4aa85555",
x"555528002aa0a9484003ffffffffffffffffffffffffffffffffffffffffc8528aaaaaa94aa15555",
x"555400a82aa0a92822a3ffffffffffffffffffffffffffffffffffffffffc852a2aaaa942aa15555",
x"55018a2aaaaaa4a8a8a3ffffffffffffffffffffffffffffffffffffffffc854a8000002aa855555",
x"54289280000002a150a3ffffffffffffffffffffffffffffffffffffffffc854aaaaaaaaaa155555",
x"522400aaaaaaaa096a93ffffffffffffffffffffffffffffffffffffffffc8552aaaaaaaa8555555",
x"52852200aaaa80845a53ffffffffffffffffffffffffffffffffffffffffc85542aaaaaa80055555",
x"52a962a100002a851543ffffffffffffffffffffffffffffffffffffffffc8550000000022a05555",
x"51a9518515450a510003ffffffffffffffffffffffffffffffffffffffffc8546a15155aa2aa1555",
x"54645046141045005503ffffffffffffffffffffffffffffffffffffffffc851aa8456aaa2aa8555",
x"5501051a114860555503ffffffffffffffffffffffffffffffffffffffffc851aa805aaaa82aa155",
x"5545552a042868555503ffffffffffffffffffffffffffffffffffffffffc851aa806aaaa80a0055",
x"5545546852a868555523ffffffffffffffffffffffffffffffffffffffffc8516a446aaaa0106a15",
x"554554a100005a155523ffffffffffffffffffffffffffffffffffffffffc85455282aaa0011aa85",
x"5515500406a05a155523ffffffffffffffffffffffffffffffffffffffffc85500a800000011aa85",
x"54550452056056855523ffffffffffffffffffffffffffffffffffffffffc85554a42a000211aa85",
x"5454544a000015455523ffffffffffffffffffffffffffffffffffffffffc85555002a0028516a45",
x"515451405aaa80055523ffffffffffffffffffffffffffffffffffffffffc8555555000a80545515",
x"4154511056aa05555523ffffffffffffffffffffffffffffffffffffffffc855555505aa28550055",
x"4154050a1568a1555523ffffffffffffffffffffffffffffffffffffffffc8555554a0006a155555",
x"4554550a4001a1555523ffffffffffffffffffffffffffffffffffffffffc8555552a5145a155555",
x"55545529155468555523ffffffffffffffffffffffffffffffffffffffffc8555552945516855555",
x"55551429055068055523ffffffffffffffffffffffffffffffffffffffffc855554a915516855555",
x"55554000115100215523ffffffffffffffffffffffffffffffffffffffffc855554a515546a15555",
x"55555155515155a15523ffffffffffffffffffffffffffffffffffffffffc855554a455545a05555",
x"554051a945505a850123ffffffffffffffffffffffffffffffffffffffffc855540a455551a10555",
x"982a0069499856806828ffffffffffffffffffffffffffffffffffffffff289982a0119990055099",
x"52aa46a9455115a1aa8a0000000000000000000000000000000000000000a1552aaa945546aa9515",
x"4aaa91a551515696aaa2aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa8554aaaa94554aaaa945",
x"2aaaa55552615556aaa800000000000000000000000000000000000000002662aaaa54664aaaaa46",
x"2aaa955551915555aaa899999999999999999999999999999999999999999992aa9551998aaaaa49",
x"40000000066400000002666666666666666666666666666666666666666666640000066660000026",
x"aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa",
x"66666666666666666666666666666666666666666666666666666666666666666666666666666666",
x"aaaa80028002a00aa00aaaaa8282a00aa00aa00282828282aaaaa002a00aa00aa82aaaaaa00aaaaa",
x"aaaa2aa82aa88aa28aa2aaaa28288aa28aa28aa828282828aaaa8aa88aa28aa2a28aaaaa8aa2aaaa",
x"aaaa828280282828a028aaaa28a82828a028282828282828aaaaa02828282828a2a2aaaa2828aaaa",
x"aaaaa28a8aa828288aa2aaaa2aa828288aa2282828282aa8aaaa8aa828282828a28aaaaa2a88aaaa",
x"aaaaa28aa02828282802aaaa2a2828282802282828282828aaaa28022aa22aa2a28aaaaa2a88aaaa",
x"aaaaa28aaa2828282828aaaa282828282828282828282828aaaa2828280a280aa28aaaaa2828aaaa",
x"aaaaa28aaa288aa28aa2aaaa28288aa28aa28aa88aa22828aaaa8aa28aa28aa28aa2aaaa8aa2aaaa",
x"aaaaa82aaa82a00aa00aaaaa8282a00aa00aa002a00a8282aaaaa00aa00aa00aa00aaaaaa00aaaaa",
x"a00aa0028282800280028282a00a8282aaaa8282a002aaaaa0028002a00a82828002a00aa00aaa82",
x"8aa28aa828282aa82aa828288aa22828aaaa28288aa8aaaa8aa82aa88aa228282aa88aa28aa2aa28",
x"2828282828a88028828228a8a28a28a8aaaa8aa22828aaaa28288028a02828a880282828a28aaa28",
x"282828282aa82aa8a28a2aa8a28a2aa8aaaaa28a8aa8aaaa28282aa88aa22aa82aa88028a28aaa28",
x"282828282a288028a28a2a28a28a2a28aaaaa28a2828aaaa2828802828022a2880288028a28aaa28",
x"2828282828288028a28a2828a28a2828aaaaa28a2828aaaa282880282828282880282828a28a8028",
x"8aa28aa828282aa8a28a28288aa22828aaaaa28a8aa8aaaa8aa82aa88aa228282aa88aa28aa22aa8",
x"a00aa00282828002a82a8282a00a8282aaaaa82aa002aaaaa0028002a00a82828002a00aa00a8002"
);

constant PAUSE_SCREEN : rom_type := (
x"aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa2a8a2a855555555555",
x"aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa288a28aa15555555555",
x"aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa80a200aa85555555555",
x"aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa8282aaa85555555555",
x"aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa80aa8aa1555555555",
x"aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa8a2aaa821555555555",
x"aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa2a0aaa2a81555555555",
x"aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa28aaaaa8aa1555555555",
x"aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa8555555555",
x"aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa8a8aaaaaaaaaaaaaa155555555",
x"aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa28aaaaaaaaaaaaa2155555555",
x"aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa2a80aa2aaaaaaaaaa8055555555",
x"aaaaaaaaaaaaaaaaaaa800000aaaaaaaaaaaaaaaaaaaaaaaaaaaa8aaa228aaaa8aaa22a055555555",
x"aaaaaaaaaaaaaaaaaa80aaaaa0aaaaaaaaaaaaaaaaaaaaaaaaaa88a28288aaa2aaa228a855555555",
x"aaaaaaaaaaaaaaaaa82aaaaaaa0aaaaaaaaaaaaaaaaaaaaaaaaaa0a8a8a2aaa88aa828a855555555",
x"aaaaaaaaaaaaaaaaa2aaaaaaaaa2aaaaaaaaaaaaaaaaaaaaaaaaa8282802aa8a02aa882855555555",
x"aaaaaaaaaaaa00000aaaa8002aa8aaaaaaaaaaaaaaaaaa2a8a2aaaaaaa22aa8a8aaa828155555555",
x"aaaaaaaaaaa0aaaaaaaaa1150aaa2aaaaa8a8aaaaaaaa288a28aaaa8aa82a88282a8aaa155555555",
x"aaaaaaaaaa0aaaaa000a845452aa2aaaaaa28aaaaaaaa80a200aaa8a2aa8aa08888a28a155555555",
x"aaaaaaaaa8aaaaa05552115444aa8aaaa2a80aa2aaaaaa8282aaaaa22aa8aaaa22a22a2155555555",
x"aaaaaaaaa2aaaa815540115144aa8aaaa8aaa228aaaaaaa80aa8aaa80a882a8a08a80a0555555555",
x"aaaaaaaa8aaaaa055540055114aaa2aa88a28288aaa2aa8a2aaa2a2aa2a0aaa20220085555555555",
x"aaaaaaaa2aaaaa1555014545152aa2aaa0a8a8a2aaa8a2a0aaa22a8aa0222aa20088015555555555",
x"aaaaaaaa2a80284555055544552aa2aaa8282802aa8a28aaaaa80a8a2808a8a84101555555555555",
x"aaaaaaa8aa2a884554055514552aa8aaa88000aaaaaa80aaaaaaa0a208222a285555555555555555",
x"aaaaaaa8a8aaa04554155511152aa8aa20a82aaa8aaaa02aaaaaa200008088085555555555555555",
x"aaaaaaa2a2aaa04550155451152aa8a28a8a2aa8a2aa28aaaa2aa882802002015555555555555555",
x"aaaaaaa2a2aaa04550555444552aa8a08aa02aaa22a2882aa28a8222a00800555555555555555555",
x"aaaaaaa2a2aaa2114055514454aaa8a822aa08a282a8808aa888a00aaa0a09555555555555555555",
x"aaaaaaa2a2aa0a1141555101542aa82aa8a28a28a8a0a22a882a202aaaaaa6555555555555555555",
x"aaaaaa8aa2a88a8401554501542aaa82a0a81220a0aa0088808a082aaaaaa9955555555555555555",
x"aaaaaa8aa8a82a8405554405548aaaa8aa28142a20280820202020aaaaaaaa555555555555555555",
x"aaaaaa8aaa282aa105551405528aaaaa2a01150a0a02020000880aaaaaaaa9955555555555555555",
x"8aaaaa0aaa80aaa11555101552a2aaaa80550540008880155228aaaa2aaaaa655555555555555555",
x"8aaaa88aaaa8aaa84554101552a2aaaa8155054054000055508a2aaa80aaaa955555555555555555",
x"0aa2a2aaaaa8aaaa115400554aa2aaaaa15505415500155542022aaa822aaa655555555555555555",
x"a228a2aaaaa2aaaa845000554828aaaaa1554541555555552080aaaa888aaa995555555555555555",
x"82888aaaaaa2aaaaa10001552148aaaaa155454155505550080aaaaa8a22aa655555555555555555",
x"a8a28aaaaaa2aaaa805001550410a02aa85545515545540080aaaaaaa2a8aa995555555555555555",
x"28022aaaaaa2aaaa1504055412848a80a8555151551402aaaaaaaaaaa800aa655555555555555555",
x"2a8a2aaaaaa2aaa8405005544a848a8a285551515410aaaaaaaaaaaaaaaaaa999995555555555555",
x"88a22aaaaaa2aaa12a0541512a848aaa285551515442aaaaaaaaaaaaaaaaaa65aa66555555555555",
x"a0282aaaaaa2aa84aaa01404aa848aaa28555150544aaaaaaaaaaaaaaaaaaa99aa99955555555555",
x"aa022aaaaaa8aa84a2028002aa84a2aa28555554540aaaaaaaaaaaaaaaaaaa65aaaa655555555555",
x"aaaa2aaaaaa8aa84a8a8aaaaa884a8a8a8555454542aaaaaaaaaaaaaaaaaa999aaaa995555555555",
x"aaaa2aaaaaa8aa84a082aaaa8284a8a2a1555454542aaaaaaaaaaaaaaaaaaa66aaaaa65555555555",
x"aaaa2aaaaaa8aa84aa88aaaa0084aa0aa1555455552aaaaaaaaaaaaaaaaaa996aaaaa99555555555",
x"aaaa2aaaaaaa2a84aa28aaaa0884aa2aa1555555152aaaaaaaaaaaaaaaaaa666aaaaaa5555555555",
x"aaaa8aaaaaaa2a84aa20aaa82a12aaaa85555555152aaaaaaaaaaaaaaaaa559aaaaaa99555555555",
x"aaaa8aaaaaaa2aa12a00aaa8aa12aaaa15555555554aaaaaaaaa2aaaaaaaa95aaaaaaa6555555555",
x"aaaa8aaaa8008aa12a00aaa8aa12aaa815555555554aaaaaaaaa80aaaaaaaa9aaaaaaa9555555555",
x"aaaaa2aa81550aa12a80aaaaa842aaaa85555555554aaaaaaaaa822aaaaaaaa6aaaaaa6555555555",
x"aaaaa2a0155542a12a80aaaaa84aaaaaa1555555554aaaaaaaaa888aaaaaaaa6aaaaaa9955555555",
x"aaaaa8a8555552a842a2aaaaa10aaaaaa8555555554aaaaaaaaa8a22aaaaaaa9aaaaaa6555555555",
x"aaaaaa0a1501440a142aaaaa842aa0aaaa155555554aaaaaaaaaa2a8aaaaaaa9aaaaaa9955555555",
x"aaaaaaa0155412a081402aa8122aa22aaa8555555552aaaaaaaaa800aaaaaaaaaaaaaa6555555555",
x"aaaaaaaa05550aaa2815400148aaa22aaa8555554552aaaaaaaaaaaaaaaaaaaaaaaa999555555555",
x"aaaaaaaa20550aaa8280155422aa8a2aaaa155554552aaaaaaaaaaaaaaaaaaaaaaaaaa6655555555",
x"aaaaaaaa28002aaa842a80028aaa8a2aaaa155554554aaaaaaaaaaaaaaaaaaaaaaaaaa9995555555",
x"aaaaaaaa21542aaaa1002aa822aa28aaaaa155555154aaaaaaaaaaaaaaaaaaaaaaaaaaaa65555555",
x"aaaaaaaa0554aaaaa0454000a2a8a8aaaaa8555551552aaaaaaaaaaaaaaaa000aaaaaaaa99555555",
x"aaaaaaaa1554aaaaa2115550a8a8aa2aaaa8551551552aaaaaaaaaaaaaaa85550aaaaaaaa6555555",
x"aaaaaaaa0550aaaaa214554028a8aa8aaaa8555554554aaaaaaaaaaaaaaa85555002aaaaa9955555",
x"aaaaaaaa0008a2aaa285151228a2aaa0aaa85515545552aaaaaaaaaaaaaa15550054aaaaaa555555",
x"aaaaaaaa8aaa22aa8aa155522880a0aa02a85515551554aaaaaaaaaaaaaa154055552aaaa9955555",
x"aaaaaaaa8aaa82a88aa8555288288a0aa8a855155515550aaaaaaaaaaaaa155555552aaaaa655555",
x"aaaaaaaa8aaaa0a80aaa154a80aa2aa0aa28554555055550002aaaaaaa00555555552aaaaa955555",
x"aaaaaaaa8aaaa2028aaa852a20aa2aaaaa285545554155555542aaaaa054555555552aaaaa655555",
x"aaaaaaaaa2aaa2aa2aaaa0aa282a8aa000a8554555405555555000000554555555552aaaaa995555",
x"aaaaaaaaa2aaa8002aaaaaaa228a800aaaa85541555015555554aaaa1551555555552aaaaa655555",
x"aaaaaaaaa8aaa8aa2aaaaaa88aa22aaaaaa855405554015555552aaa1540555555550aaaaa995555",
x"aaaaaaaaa8aaa8aa0aaaaaa8aaa0aaaaaaa8552a0015000005554aaa15400555555002aaaa655555",
x"aaaa8000002aa8aa00aaaaa2aaa2aaaaaaa1552a2a81502aa05552a815440015550004aaa9995555",
x"aa001555554aa8aa0a02aaa0aa8aaaaaaaa15528aaa8552aaa0556a8155100000000050026655555",
x"005555555552a8aa20a80008aa2aaaaaaa8554a8aaaa154aaaaaaaa8155540000000454a80005555",
x"555555555554a2aa28028a0228aaaaaaaa1556a8aaaa054aaaaaaaa80555540000054552aaaa0015",
x"55555555555522aa28a80028828aaaaaa8556aaa2aaa2a02aaaaaaaa0155555001551554aaaaaa80",
x"55555555555542a8a2aaaaaa282aaaaa82aaaaaa82a8a8a8aa8000000055555555555554aaaaaaaa",
x"5555555555555428a2aaaaaa0282aaa82aaaaaaaa802a8a80000aaaa0015555555555554aaaaaaaa",
x"555555555555554000000000aaa80002aaaaaaaaaaaaa800002a8000a001555555555554aaaaaaaa",
x"555555559999999999999999aaaaaaaaaaaaaaaaaaaa000002a02aaa0800055555555552aaaaaaaa",
x"5555555555555556666666aaaaaaaaaaaaaaaaaaaaa800002a0aaaa8a20000155555554aaaaaaaaa",
x"5555555555559999999aaaaaaaaaaaaaaaaaaaaaaaa80000a0aaa8aa288000000555402aaaaaaaaa",
x"55555555556666666aaaaaaaaaaaaaaaaaaaaaaaaaa000028aaaaa2a8a200000000002aaaaaaaaaa",
x"555555555555999999aaaaaaaaaaaaaaaaaaaaaaaaa0000a2aa2aa8aa220000000002aaaaaaaaaaa",
x"5555555566666666666aaaaaaaaaaaaaaaaaaaaaaa000028aaa8aaa2a288a0000aaaaaaaaaaaaaaa",
x"55555555555555599999aaaaaaaaaaaaaaaaaaaaa0000022a2aa2aa80a8a2aaaaaaaaaaaaaaaaaaa",
x"555555555556666666aaaaaaaaaaaaaaaaaaaaaa800000a2a8aa8aaaaaa22aaaaaaaaaaaaaaaaaaa",
x"55555555555555559999999999999999aaaaaaaa000aa0a2aa2a8aaaaaa22aaaaaaaaaaaaaaaaaaa",
x"555555555555555555555556666666aaaaaaaaaa002a88a2aa802aaa000a8aaaaaaaaaaaaaaaaaaa",
x"555555555555555555559999999aaaaaaaaaaaaa002a22a2aaaaaa00aaaa8aaaaaaaaaaaaaaaaaaa",
x"5555555555555555556666666aaaaaaaaaaaaaaa002a22a2aaaaa0aaaaaa8aaaaaaaaaaaaaaaaaaa",
x"55555555555555555555999999aaaaaaaaaaaaaa002a22a8aaaa0aaaaaaa8aaaaaaaaaaaaaaaaaaa",
x"555555555555555566666666666aaaaaaaaaaaaa002a82aa2aa8aaaaaaaa8aaaaaaaaaaaaaaaaaaa",
x"5555555555555555555555599999aaaaaaaaaaaa000aa2aa8aa2aaaaaaaa8aaaaaaaaaaaaaaaaaaa",
x"55555555555555555556666666aaaaaaaaaaaaaa000000aaa00aaaaaaaaa2aaaaaaaaaaaaaaaaaaa",
x"55559999999999999aaaaaaaaaaaaaaaaaaaaaaa800000aaaaaaaaaaaaa800002aaaaaaaaaaaaaaa",
x"5555555555566666aaaaaaaaaaaaaaaaaaaaaaaaa000002aaaaaaaaaa8002a81400aaaaaaaaaaaaa",
x"55555555999999999aaaaaaaaaaaaaaaaaaaaaaaaa00002aaaaaaaaa821002a84552aaaaaaaaaaaa",
x"5555556666666666666aaaaaaaaaaaaaaaaaaaaaaaaa000aaaaaaaaa2842a02a1550aaaaaaaaaaaa",
x"55555555999999999999aaaaaaaaaaaaaaaaaaaaaaaa0002aaaaaaa8a12aaa801554aaaaaaaaaaaa",
x"5555666666666aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa8002aaaaaaa084a800010554aaaaaaaaaaaa",
x"555555555559999999aaaaaaaaaaaaaaaaaaaaaaaaaa8000aaaaaa04128202005052aaaa80aaaaaa",
x"55555556666666666aaaaaaaaaaaaaaaaaaaaaaaaaaaa0002aaaa8844a0aaa80550aaaaa112aaaaa",
x"999999999aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa0000aaaa2844802800014aaaaa8454aaaaa",
x"55566666aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa80000aa8a8120002aa812aaaaa1454aaaaa",
x"999999999aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa0000002a810002aaaa0aaaaa85154aaaaa",
x"66666666666aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa00000aa84100aaaaa2aaaaa85154aaaaa",
x"999999999999aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa80014aa04542aaaaa2aaaaa14554aaaaa",
x"66666aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000015281154aaaaaa02aaaa14554aaaaa",
x"5559999999aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa8000545405152aaaaaa282aa854554aaaaa",
x"666666666aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000155544514aaaaaa8aa802851554aaaaa",
x"99999999aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000155545452a02aaa0aa854051550aaaaa",
x"666666aaaaaa8000a00a0202a02aa002aaaaaaaaaaaaa0001554154408a8aa02aa155151552aaaaa",
x"999aaaaaaaaa800080020202800a8002aaaaaaaaaaaaa0001554500000aa00002a154151552aaaaa",
x"6aaaaaaaaaaa800080820202800a0202aaaaaaaaaaaaa0001514454000aa80000215455154aaaaaa",
x"99aaaaaaaaaaaa808082020200020202aaaaaaaaaaaaa0000501455140aa80000015555150aaaaaa",
x"666aaaaaaaaaaa808082020202020202aaaaaaaaaaaaa8000055455450aa80000015555102aaaaaa",
x"9999aaaaaaaaaa80aa02020202020202aaaaaaaaaaaaaa0005554555142a8000001555504aaaaaaa",
x"66aaaaaaaaaaa000a002020202020202aaaaaaaaaaaaaa8005554555452a8000000555454aaaaaaa",
x"99999999aaaaa000800a020200028002aaaaaaaaaaaaaa800155455551408a00000015454aaaaaaa",
x"666666aaaaaaaa8080aa02020002a002aaaaaaaaaaaaaaa00000015551450aa0000005452aaaaaaa",
x"999aaaaaaaaaaa80820202020002aa02aaaaaaaaaaaaaaa80000015554514aa8000001442aaaaaaa",
x"6aaaaaaaaaaaaa80820202020202aa02aaaaaaaaaaaaaaaa00000055545152a000000000aaaaaaaa",
x"99aaaaaaaaaa8000820202020202aa02aaaaaaaaaaaaaaaa800000555515548000000002aaaaaaaa",
x"666aaaaaaaaa8000800200020202aa02aaaaaaaaaaaaaaaaa8000015551554800000002aaaaaaaaa",
x"9999aaaaaaaa8000a00a800a0202aa02aaaaaaaaaaaaaaaaaaa80005554512a80000aaaaaaaaaaaa",
x"66aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa0001554542aaaaaaaaaaaaaaaaaa",
x"999999999aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000014054aaaaaaaaaaaaaaaaaaa",
x"55566666aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa800001514aaaaaaaaaaaaaaaaaaa",
x"999999999aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa00005544aaaaaaaaaaaaaaaaaaa",
x"66666666666aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000005550aaaaaaaaaaaaaaaaaaa",
x"999999999999aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa000001550aaaaaaaaaaaaaaaaaaa",
x"66666aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa800000542aaaaaaaaaaaaaaaaaaa",
x"5559999999aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa8000002aaaaaaaaaaaaaaaaaaaa",
x"666666666aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa002aaaaaaaaaaaaaaaaaaaaaa",
x"55559999999999999999aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa",
x"555555555556666666aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa",
x"555555559999999aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa",
x"5555556666666aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa",
x"55555555999999aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa",
x"555566666666666aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa",
x"5555555555599999aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa",
x"55555556666666aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa"
);

-- Begin Behavioral
begin

SetColors : process (Clk, Addr)
begin
    if falling_edge(Clk) then
        TitleHorizontalColors <= TITLE_SCREEN(to_integer(unsigned(Addr)));
        PauseHorizontalColors <= PAUSE_SCREEN(to_integer(unsigned(Addr)));
    end if;
end process;

end Behavioral;


