��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�ϗ7�#���H�����u�g[iˬ���t|�3���ҥ�ys�B�@Yq�"F}�\"QY����#�ڇ7�\ӷ��繟��1W�k���q�u ���{�m)RM�S|@�����ͣz��yʿG��O�Yg>�s$h_!��-~���=wx�=�M�����/�mb�K#�� ��1��W�i�{,?�EM�N�0�K
䧣�:39ok^�(��-���V�f���Sk�	����}ؖŸ�*����~������6l@ޱ����t����_.��±7�Eۨ[�ܐb\T�8�����"��!'���^C�he�K�Zw��J�;��E���a�BnB��lje8�i�U��^w�K�@ܚ��^<'�������������a}��a��W��S��!�P�:�ޓ��|=ǎO�k�σf&�_ K(yǦ�+F{v5�X�x!}e�y�D��"љn3]��6:�Ѳ=&:_��h�,�klf�es�4�=|��-�#3��r�E8m>�e7�{�~w���O3��{	 X�n���7��[��{d�mҫFG�6�ݝZ���4́���GF��yw�D��Օ��挹O����[�K6���L���ڹ�\Z'�
���lS}d}��w7�� ^$�j_��묡X<P�`��&X���xRq�y��G���R��B�}[�b50t��j�k\��Ju�a�V�ؒ���w�\%RF�Z�購�:*EO�GT+���,��B�/�9K�5J���t	���y"q��yǕR�<�]���>{�t�f�'z�(*��l�����'J|N�]�F����Yz�ȅy��/��)�B��
�vu`o9M5|�Z�e������gM"���C�W��f,�o�`��<��Xk�:�s#�T��/q�PC���k�!}5������j��b%׊a1-�b��\%猢��S������Ew�Z���UYwds�i��;�IT'q��z9}j��!/m�n��4�Z������ء�\��0d��>�fZ{�>�Q���}o�x�/=̪Y�I�s<T�y-���G���_�җ���2���5�g�$K�+�'y��wj�%��� ����s�ٸe�p{��V�$C����FQTX5��)w�"��c��Lg+Z�fvV@4�ZP�>l���
�U��������tAĪj�k��V����>lv�C�/8��M�jR0�:q����Tԅg%�L�:�����t}W�/vF�XȰu���*_=�Ҧ�/W �W�J��k2|�v����Q�o�2�l� �@��n�S&E����q;�Ǹ�(�b�?��&�pAM�� k;Eb���7��U�U�k�и}8�+9$��'����ݧa#{�~P�C@�u`�#����]�S�N{"C=l
�i��+*<�L�n�k��STA��s�%�X;�y��@����L����n��e���-�4���=���t�X�	���B�`�K�C���Ɍb��8!5te���i� �������9�E�y�w��ܺZz�
�5�_�w�.W%x���|�	
�Z�� /��x���f�-H>��|�)O�(�x��:E��&��Ͳ�Q����<>�E������B����
\�t΍��9��Ȟ��\���$�z`�� �1n@4/��e�P��$���u-��?�J�$?���Q�Mʕ��[��y��ن@0ha,��t�H���OD0�p�{O��M=f~-�G����(*��!m�Es'�#�A~�G���yk"�ї�����!A.���Qձ�&Yeis?ޖ`r4��9��7H�͚J9i�Ň�yʣ]��,�y��)�Wz1����?����Wt����� ���� �mT��"�\<��o�����D���^ϝe�x鞾�F̂���ˁ��ͪ΢:yz���Jc
��CN�!=�,�]$a�����Ù���2���rTc���Z�=HZ�$�Z��^T�{)�ȧ���_ׇ߹k ݧ �dظ�z����*����D��٥=ɬWb�	օ�����^���Ar�pLPH�7��G(�.O�]\��Snf�ǯy��(za:e�^������.�Ƭ�r}�GMP�s �Ǭ�����O�x����Y�T��3��`��3h�s:����\2�d�;n-�q8���FW��>3�|o�
|�ÿ��F4I����[Lb�8��9'�Yj�l���[T��i�V��p���eƤ��h�9���`=����[Pf��c���#����4�7����Y.@�ݧ��{��Q�MDm��D������C��2��]�4���vK��B����s�6'.s;�Z�U�e9J�:9�7��@T�_��ꐜ�M�x��>�`�� ���"�k�(V�я�����5��GS����ׂk�M���I	ǳS��Q�N��P�ĜF�GA���Wy�j-���D�k�*��M����ՒJ	�q���Y۩>q�S���R�(Em�F��\���-�h���Pj	M4oı����DN�����(,�,�|��SO!A�5��.��2�ɉz�	�K���q�'�=[ʭ|LX��Q�h;vn�S;̝�Є�%/o�f?*���[�B*�z��K4��)�D�gz��+.ݕ��c��%�V{X,,7+M�0cc��;L�W���zo��ϖQ���"�L7�k��1�鲾ě@�uo#]��` �00�v�3)��e�o�g9Д�(�e�$��5�z�m�7*'��
�.�J��ly�L:,ۨWu0B٤����?��RĘB+%yY�|�Q@������¯C>�<卓���<X�dI���I:�!�r�4+#(lpؒ&1���эb_�+V"������a!!�h4�B��PS@ {4�i.����eG�\�w9v��<��pp풥�OYY�0������Co�gFFp�[�|o�s��u��-W/�Hx�o3p�+F�;Lг6]6b��$�^W(�,ބ$���(�?�g&kyt_�e���s5���VE����{l8ݎ��Z�x�'8�^+��Wl8˧N�]v�Xѡ�t �m\K ���a����)\�$J{�[�=�4��h�}�iy2Z��TDy2@��k�N0��~���qt�x)�{��N<��LW`��uT�*���(�;�)��)���@N{��'zoT)G� B|e�eH\�(8���@�,�V�6����r��_8K�E:��&w �aeC�&f.f\*������2�e��C����<���
0�?��u\kYA^M��*��i^�X	��0]Zs��))�z	��l��8k�aNe2��i��3V5��]��zv��� f�\��$��Oƺ����Ni.�q-�Ӭ#��X�	O6�<�)��c�Xͱ�3��X�Qw���8RJ�x�(��xsC�-�
;Տ����px��'lHR
��Z��{|�{�1,
 �e7ų��	f��������~�GPV�S5U��0���(�ẗx4��������W��H;�*����j�;��������f�������D�Q�H�Nڡ��gT�Aw75��7�:�C�X��4�>�<%�i�Z;n5�VJU}!�0��zu3���ky��`0��M��
��j����eqw��T�xvB�c�1EzhMP]0X�X
"4p@HHW$�ik\9��D�{����i��Ԉ<�2M�v���,�@-q�%v2���,�=��埱�lѕ#��
%Z˓u��O�
�q�:0m����K�Pu�!0�;���j�\�Kyv�k[�0z�GN����ժ��R�Y8-&����i�]d���� ǹҷ��c�&�qO�&o.F�Eg�=A#%0`�Jn��U5�I!�d�l�J�J���V2Ylie�K��:_BĘ���;�����.B�|d��`�g�- {�y�Jl��L��&r�6 x�M"�p{�[�{Wc�=�!�ٓ.ۓۋ_��I[n^�� L^�
��2���I�R@쒬���H�n}��ఉ�y�fÅ	���>�,r�-�-^�<1�L��$��h˰���L��X�ibI/�K�J��jXc�n��w<�A�J��ȅ?����N�ݤ�z��5H���ߺ�=x��S�ˉVH�x���Ր����p��O(#	�ӽݸ�� '���⩊<0�v�o����V*��Kr-�I
�w		Ŗ��i��|����9|��N�3�
(=��0Sh�@˔��f��Un�6�V5Վx����o��B<�99?P.��/ H����gY#0�<	��� ��+PZ�E�V��)�J
��s���.�N�ΙyŽV���_I��O,��`�'��<|��YЗ�[�QҨZe�T��B�0\�R�:�&�>�B�Nݠ�,ʝ����/��� u�=A����#��d�
z�U�x�5����T��4�sK���m��E5�rfcg9bx���ʶN��V!�Y������)#-D�+)��9D�$���+iV�9�SaP�	�p�~>r�o���n17�7RRZA77e�)*D���˄ߣ�d�f��������)�%��< J�v��)4nO�D�Q�)�wDX5�@a��=�;�7��a_w�OR�zw�r睟�;1�?���17�0F4OaQ���܎��Fk��bp�k��o{��u�������?z��dl�+�H[m��5��xg�#3&4}����J4�
(U��Q�-���3x�T&4H��(����|"��Z.��
���hN���Llk~n�q�A��1��x��Gޓ����bt$���pԸ�P��K4Ķp����w�Kf,8{k�dA�i�p7��֩�i�~}�G�d�Jn/��1?>�n,�i~�n�sh��D���g)O5X��u$+�f���V�z���\(xL՝\�GaIrE/`;�&���m.�7
�\��y4�Ie^S��/u���V1���?���B�e[ '��{��SB� *6���k��� KR����z�����h��g�x�ǭ�ʧ�Č����J;)s'W=w���z�9Ich)=�_�#8�{���\����=�/�`/����ԂapQ�����X�+�^j���`0H�t^͋�Z���u�R�Nl)$�^�w�*<�xG����.����Y���Qp�wu�y`����R�Zj��@�ery���y��	ܠ���w���$�]u`1�f���pd]ӏj��u��&�fU��¤��7��K�>^FA@gp�
��J��N�l��[P��k�Q�����Fy���Un#g	��g��'�mO*��P���N���1�>W��c��l����Nֈ�=��k���6�fsm;�\o��m$hjAW~$��a��o��`�@�c�=7»9u�{^��%�ؤv�F|{c�;ǉ+ac B�f�R�3�g�S��J�Z8�)р���F�OA'y�[��⫖%
�L �0�}żА�f���,^���kи�>l���Hf����j��G%�=�ܣr����dYD}q �y��Hf�
x����F���8#�B�R����s�[�m�Ow�C��"���F)�ޜ6iP��k��ӹ�z����T�;�o�Q���×HE���n� ���z�f��?:N�s��(�j��W*s��u�f8}�U�K5�#a�5+��V�bKI�R�K�rQ�a|�U]��xq�����n���]&%�\�/�a^�:�3Jkc�'l�n��ǎ�5(0Hש-�u��J�z{���@�1Wӆ�̀��������VCQ	K%kl�b.�<�Sx����c�Ü�B�w�1ڙb;u��Ʊ�������50X�hr2�G:�����JI�'�IO�V;Q)+�V���.��wh��.4*�gH:	�(7-��[X�DT�L���j,ӏ[���e8�'xd�O���*���Yrnx(������x&,K�<���d�SU�ߗ��J	�7��J?H�ڒ�@�f�p�"ћT�#%�E/}�K����>:E�����k�R.��Q/��7���%�ʪ�b��|�/1�b���谕�TS���~���*�5GKf�/qk����F��TkF'��ReY�KmVv/����-B2 �`��j$����M�FGC�`Y����EB�I�e����P]N/:��9�_�����N.��s��s���4]�aI�5�
�l��N�M��5����W�!�]f[���h1Ħ	��Ń�_ZX�l�է賁�U^Y�E2|��lƉ��^[)�G�����8�%2�0X�D�t��¿?B�O�7���ū̠�8�N�"8�;-�j!����Wk�}/����ȳr�6�(�e�}T��2�U�P+@ސ�ӆ���AϮ�R7D�D�/+��oC�1�U�#�i��_p�4�3��G%�]#��NwN�zY��Vۧth���������TL�`�3g�;�e�a�@L?���t�mOWX�p�s:�V����a�����C�!_�I�w�)���a�������xُ�+����R ��(T�ierUc�4���t+!��cO0=n��+�CDp�!}g0��I���jH �A;:.4bYv��#�w�O���c9�@	�K�5���Z��
�$.��c�+���cr�3d��$Ч��ˬ$�G�-��n�%L������Fdi2������t�H�y�,���v �$�=Ͻ���9��[��r��5��9�J>��T,��X����ʟ��EQ��)|,��C�]8�����y|dާ*��D~����#Un+~.�$�x#b��v4����v�=�Ohيr_���1敾W�	������p��1�t�.4æ�e4~��"8/V������|*������贼�((@��]{Z��H�� ���\�s�w�G���q't����[!`t,wNV�8㾽�-_q3��hD�6H���%fv-��4���a8��5�N:�)�[���_l��F�yXX�������+��x&`,��Z�`��7?g�/b�ɀ �9����/���o.1Ʒv4k=��z����Xn���0�Y�4!���A�!���mK�{��FE��Ww8��qeVd(�%J¹���0��ܹ��;L#0ݱ=���]P�j��"]��i�CC�&�GZ�VY�+#C�a�@E@���2�� -"'�xf��s��6�mY2.	��P/�G��$s|��AU.�M=��+p«3TF�Y�@t,�Qb
��5�Xj|�*8��n4�]��ii�l��Y6,c��1\���&�����k���e1�m�<������T�=:�#��Uy:2�� a�C6�0�gܛ�q,Ix����Z����-�e�JB� jnJ`��~�1�q��ڀ���2�j�Q:�@?b��1��;��,x&b '�8?�`S#��B����&��iB�]@�L�#�/o[�oI�
�:�4��o�ͬ)�K���@��
Nf<$���m/!�"�׏��3� �����T��Ƒ��=��y�-�r�1! ��1ix_����v�3BR7���I�]��)PS�ҧ��f_kA����Q?m�������hc���P�z%��,~k���w�Ͷ��Ξa�Q��ܪr/�t�EuP���6�f�������a�����W_�J@KL�9�`�#��-疩/bl�FW!1�����*�����wZ�)��f���ԃ��J�A�.�h�@C'�����*�T�~��"=��rL' �vC���I�{�- ���&!K(�.�s�����P-��4�Fo���E��w�s� ⢽]���-\O'�߹d�U�	�jH��ԝf4�;rG*D�_6������~P!Z?�;wА�T�T8]�_�>�)M�����tXz=�{���4��rץ(i]�v��Lhϟ�fś!Y�K��m#�/���~�J�	����*�o#\�H�!>3}-����Nl��M�m�__o�`���R�5���R�e���'5Q�Yo����Ø��ԡH��U��t2�o�	�		�*��c�lxe �WEmK��z2��347Ԛi���䩰��bl�Y~��f��Wؾs�ڝ�&Ϳ�	���~'k�gC'���&7K� ���œ9!�;�Ш�"�9����SrEƷ�������Wo0�f%l"�A�M������Nx�9�~#�-Oy�e������Yʛ�=P�[\�o���)ga.�� C��߶gk	w\���w9~l��z5Y�ڻ(�`��,�U����<����kd<"�Fk����i 2�*߻�����m�i����*`��Zɕ��:+�5R/�,M�lb�O��.�� �s��ۓ�e���sY�j�w�P�ku�bm�D|�G'���I�;{���n��&�&��{��4fk+�[���0#��u��%�YǷ���D���ޜꤲ\yjK��~Ɯ��1l���
������i49��\odf��'����$�ۤH;�R���}	]G���T��uZZ�{@ߒOzQ�TY����!�z����ī�jL�n��m����4�sEu�Q�-�	�,5ёZ��C�*uɇ��?'�G�;Ek���ʣ�[��f�;l*�д�#�斡�{��߂��=���"�z��KR��r8]��D7X(�ﴥ��"K��$��|Ao&��v�����75jV,Nh\dΞ�� �I�%h-��C���Yy�1q*j���qN��~������]gG�L�m"k>�����:\���٦' �O\����E���׊���;��;^&ժ�k�P@�·3�z�eȲ-�N \�|�}"�h�e0�����'M�`�x�R�U�"��6�ܳ��ou�ȋ%C��������I�<R��������N�@��J�ٶ�٬�u>;����x��ýCۦ�25�N�S6� �dS�b�y������c���U>Y[|����W�D�;c)f���YY��ELtN]�wg]���.T�c }�f��$tեn�����Y?W�NO��8�w+~]_�*���2�x�e�bq���F��	��bp�$��=5-譖I-3��Bj�?"!�v���A�Q��	��%��c{>o��!�Vޤ����j����b`�P�w}� �dJs)׍Ci�Ej��$��wk���\�
����.8ɲTݑ�^�h��L��?�F��a.dZZ�d�f'gF�7d^ h�ۈ0�I�汓�=�|��^kla+�O���N
�+�S�>zxM��d��U�P��{C�L�Bv�v4̿����q���\��k�G\)/ Q砷D�ǌ}��I���1�&�����ZtN�*�H>d	�3l�V�@��`]����Q��YU��1�#K��?N&�=5��|��ž�%1&���u�)�T�ڞ��p}8��o�����y#�)�����5�5:�'�ũQי&�'��5h��{ֈ��|Q��8
�i �'Om��CK�w��=Vlos�n���a4H&+ؕ�n�{g�|VW�W���LÌ\�Ne%΄�X��h/b-�k	�joz�.�Sn�k��!Ƭ��6���Z����5�;��x@�~Q�˙�ɿ%��='�3�{#���{jᚱ���r�f`��_��+5�&Q����� +M�/���g�@�񡰧�Q�̽U��ꜿC���;��T]�a%S����y�e�e����5:	����b�m�.��Z�5�;;�a��EZE�o�N� iީt�������V^7d�pr���Rʉ5�R����W�5C	�R�y�y<(�wH�o?����.�Qp�DK�}&HG��38\h��/o�\��w<h���Dd;_�cїlX��D�^$/�ۭ̐ߠ��E��?��j�Yz��OE¡՟!U��@S}�G4zj�m=tr��0����ۼ H
�hՄ�OZM��B+���S�(��<��E��>�J�5D�k�0otN�T��Q��Gh�6���^ѷ����3��p#j/�O���� 7���n؈QXܢ���w�u��c�AX�^O~��'^�I3h]�����4sώL!Vr�7��	�g<8a���$i;�
�{0�p*�}�vv��#q�9y}֎6b���l'�Ә�D�Y�EfX�@������5p�����s~�������c�?�4��Y����?��*�s�PK2 �x���x���w��)���X��\��f��K��""�Cx���y�$~�BRvݧY������*�xUhnrY*��Z�U!�%X{�
��T�F�H^툉��s�
ncX�춼�7��\��w�v��$�T�)��w����yp����ICXuu��H�f�:�ִ���<�*Ӭ����9���
���B�ž _�ݥ����HH(C^�#-;��KZ�%�ǐ�D>���?���-9�9<Ԥ��u����_��E�[ꇘa5/Ia�f ����"z^��}H�`첒-�k�)�u:٬9�8U�6�ݎ�~A�E���D��z�h���S��b�W���A��n����*A�%�sf^ �2+�{�by��uַ�#xt�~���*� eT����N�d�����ms��+c���
[�*q�s�*��d,�b�M����͕��7�h���e���{=#�����]��0�I�q8n��h<�P����Q�O���,@4/lS�PZ�ar�&����ƕ�X�=��-P<����&�c^��d��;�`��Ve�^�5����'"'؅�X)(S&�z���J��<�vT��`�'�q�Q�a��%��6Ϳx0��hȡ�pO *u�-��Q��	?C����u����E�C���O{R>�;�Vo��]�J�~��5�:f~. ��r��ͥ|s��9T#A�g����.�����~r������96�7SROT��R��g ��KԞw���G7ߣ�6�u�tn:&��6��|l����K"�(�&�|� K�'���{|f���-ؚWy!��8��?۹�K�\�U���b	��v
�l�������WWh���x�H�����es��b���#!{%����*�-}�{NwK��RۿiX/�Z͜p1�o��nma��-0���;+��t�a�j��4Մ��i4�i��X�rp"���W����S��d椗���%�?�g/�9�c�p��x�4�w
�7@Gpr�P������o��epvRK���J��Ҥ?r����''x+s	|m��;�v���> ���IYH겆���6k���L�O���3 �^a�%y��P��+;��u��yg�`��+k\�������p�=*y�j��r�
��C#�<�^r����V�dv�r��X����!����сj-�[���.�./��T���;^����/A���0�r����3����q#��e+��V��E�L��~� ��h���}��H�]{&k>*��l0�Ne#�b�)�ҕ�8	A]�{썌��*�ʠ<�.K�fVe�fS��*63�5Ӟy�4��?�R�9ǟj�1��_���Cb ���PF4��@T8�e�����1߲H��W��gY{���)�����і+ח�lgk2�������6wq���)��v.����Y��Q� �>	�&q�`�����S������g�e��&����&6^ོ���ir�.(����r6uJbF��\oGo�
�bE1P��/�;M��6-a|�A��T�('Q!
�T�v-�S!�̈́_�9��b9->oM|c"�Y\Tn����df��+�*����-�:ni��jM�7座_��B�^�u"ͩ ��%4�s�I�s�z������z��c[�4��˦��7����+�`���S���#g�~�`�@:�s1�g2�p���[���k�$�V�ɲ+x<h&�#��fp2�A�A�7]����Y�W/%G�I�1W
��\�s.�Tu�t~kdW��~�-����Mh����=ܟl��QV�51�SX�,�]�fHWU9�h���oa�՚ ���
J��t�!�;H��~}i7�<�t�0c%D�>��q&;x�F�d�f�n�
�w�Iȯ��i7D�R� 3�p&�%��F�m>�E+n��FI�eϒ��GT�8F]?�e���rV�"�6I�W'ĉ�&dMP�B�5���5��:~��A�=j�2F�(Ø-�կ�?�|e�#2��W�nE���I���C���Q,�oe�շ�)b�!B^�h�km���L���(>���Nk��ۉ�b�Z�/e�TE2�Ͳe��6`dv8��k�����Q��j��Ks�E��q�W�Uc�"�XYz�w%%#쬏6Tx�����
���L�� $��>�;�ѻ�������ϧoe*���S�"�ǩ�E��y�8$
P7!,�E�����
�!+�Q9�c�*�@o�D�L�߫Q�Es�M���<�n��7�F�t��A0kI�Pg5����0!ͦp~i1�lՉ��C� !w< �� �}�����o���v�ҏC(;������`4wϪ^��An��m0�� �=?:1���e�-�9�mՄ�CL��g�e9�>Bv/82,�xgS	���@ ��Ly�,�����;�L'bzϦn!�g�wG^�f,c�N�/��	��N<@�k�.s�\���B�~�7�)c�GM6J�qW�]j޽�Y��Vn�ږη=yL����o�]�S6ĺX��c/a���(��.�t]т�_P�G�<c]��/�L� ?�����"���N�upwMٔ+	��fD��N��e�L˥m.��`�9Z�۰C42�_
J��B/��v�XU��L����^r�uv�r֪�-Z��v4����)r�ۣ�:4�����?\��eD�6"�4�̠-�����!V�Ug��y�9r�ujpXϽ��a�sP.h�JS��T�]��B��v�r�.ѕ?��m�'O��j�S9̌v���4������6�X�8׌��H�"p6yYF�q<�����Oׄ+��nZo��h�!�[.��b�E����`E��K6��n(N�n튱���2�P���c�'��������V n�
�]>�e��˓����O���fP�nN�Vgc���w���h�QBm�W�N��T�Z�wCX�����W�#I��W�Z�i���^�,.W��(A�C�*A�,#�>aϵa!�L>ۅG;f�=+*(����]����ϫRV�Ƭ�Ǟq{�gY�������<! d���+3�>��[�)m?��N��z�QLZ[[(M��w�ʱ�\�6�b"�޹|1Ȼ���FV���T�DID�p$+aoc�P:�t͉n�����a� 2�G�ż�����O9�=��I���T�1�S�Žp���rZ�0Q��NK7�2���N��vD�ێ�z��$2z�T�F�b��@�@o�;�I]��y���=�3�_������yd~;"�<����Y��P z�b��8Y��l7>���ϧ{�(+�q�Y/~Xt����$�.��{Ǌ۲F��m�4%Ѯ�����*	@U�"���?j֞Y�+V;|��VH���T���d*���S~k����_>��������#e�	wC_1�&�ў�!���~͹���[�k��2h��{h�UwW�>|:0�nȈ�FGe͒�%��'�����e|����b�]F7�Np,r����5Fd�!2|?�����`�i>VMT��X1)E�������p�c��*��\rfݽ�c�QsmY��J6	�q�׋V�fK%r���h��ћ���ޣI;�b@A�S+�Rqb����o_"C�������W�J�/����59t��Gd������b�<&�9�ߤ�$�N��5Z}�����U���W1�ӽ.~�3
?t"���H����T�s|��Y6�d�����N�q���bN����D��ŖL%��b���>�T�ٽ�4%<C�>W��f��`s#^���@I��dl-|�׼��0��&��K=*�G�C�kX��T2�k�RMI��Z|�����ݍ�j����6T3�����^f�p� ����~�U���:7;�f�S'ep��^�N�D�Bs�����k��%d�laB��O���*�����x㚶�wbj~�G7a���� ��)I�?,?3р�%U(M���%��6��!$e�"�:sUX;^2=�x�h��frș�����>	e�~]�U�1���\�:�2R���A;]�%�*o��:���N��Zy�T�����`�=?���Sq��JW�O		{�- w/#�S�H�P��/C����?R3|���й�zmO[똿dkfS�!�޳<g�V�a����t�N�V-� �eȪX%b�(�)#DoN}T�xNW��52Ӭ�܉�J�-���3��'���r]�DyGC&�����n��Hk�9O�[��#�����̣�%�w�C�+x�pi>S�ȑ����������~�'��+��Cv�m��IX�)n��R�"����Ƶ�S���)]G����[����IF��Ѿ
L̺�Ke�J��,�i�APV������K����a����D}h����S0EAKTCK�]��j��?�sd��A<C	åCW���NE��6	aΛ���./>��k񊯚p���&�?G�sO!,>W{��v��w=��ZJSz!*3��1*��Q���҃�0�ڐQ��m�Hΐ�3-�Mx��\�G�eQy~��#X�4ϟV��%YH�7a�0�7P�\`Q?��5V<E�*�xН��r�Z��[9nv��Z�Fb���e��8�hd�����+;:P��	�'�O����J/�e����ޮP��w�t>��k��	�����=��ɞ�*��H;`��Ǹ�*J���b�*0ko�7�W0^քىSKVzה+n�����F��tk�wh�e)Δ�m��ʝ
�Vv�k	�����
R�*3\<jm�P �pX�l��m�bڪ��J��^��������6wq��:"�TQ��(k��A�m�VlD�o�7g9�Ri.kD�����Q HdP�/p�Gw�PXTEB�&��/�dGCn�������u
�63��T��� �����{�f !;t���g������R�8�6�a��k����]��ܭѴN2�gt�6A?��YK-�$���@^}<��m9(��#�����cy!$o5:DC�ev�B����F0�'�s�1HG�	1o���Г�X����r��>��.�IPY���5�� ΃�8�\�A
��0:������_mbE�nM?C�J
����Dm��e7sAs��s�sfR]�!���F/�C�8�ܻ��)ҝ�?�s[C��x��TvBN�+.�J�ǋ��n��nkK;L,,�{L�i�i\}pB�T�B�S�}���-�M�*����0��#:�j˕! @��Me@�	9w3��`�a��ޯ���B#ߴoҵ�b~������Z� F,�ŅҾ��Ē����q��kJ���_�)��Vv�ת?
_t=�2t�1OoH��'(+l��^��`+��7��RΈ�0��7&U�o_?��'?�v�0���\O�!�<raa����n��"�_8�c�Ժ�u%~;��Q���kD��K�%V��E��^��_�W-��:lUđ���3,T{�V�Ou^/YK�x�gD��d��"3�HMkX�?�|��äje�=��;9��;��h#�f4���k�u(e���h����g�ȍ~�����e����᳸�hS�0�L�Ӵ
�R_��PE�b4�C{�99�ky*ɮ3��*���±�K���7�G�dv6��>��ہ�l�'�_cҌ�� 60��ZR�@n�j�m���꼙9+�5�*��E�h�'.�CC�6��f�|1�Ǒسp�oȬOL�N����.%�Fn�j�=cs����[���S܇��S��
��v����|��o:4i�
�X�<g],�{)�G�!��g�uV�3�ѩk���ٍ���D��]j���ғ
xL��;#�i}NxR߳��*5:I�Ȫ���� n1��gy�7��FW�tԩ�AՁ�wh�ěҬ� �"\k��#o��]���"��UP�3a]�,�ү�}@�I��RJ<�#�1����� ����դ�@o1#߻����ܠ�h}�o���3>�r�ks<�G�r��<�@�	#���
�����D�J�򘩴h�6��'��ȏ�sе��_Ri��%c�(��K�O"*AR3ϕ���)1�L z��l��~�Fu?���@Y I��<ʄ�a�'�͐����1@�|;���gw}�����X�7��)��1�9|�u\���-�4�^���	�A��]��m���l\�Nc�A�Ãg���uk��8⿈=��>�� �ܟ!EM���j����K�,��ߕ��"�,4��3�o, 3k���b諽sN�E~$6���>�b{��lɞ�����`��Z,���gB%�&lX���� ���E.��覸�ߘ_�e?&�]�� E�pS�˿Q#䔬���WUX!]�v���LIw&�,�7�u����ͯzU��6��Ȓ�[�'REd�\5Д�dϨH�H��, d7Rf�>�c�7�<o�\$<0ܪ���_9�h�q�IA�Y��*��o�l��eB�M�?̅���c4�D��PE��x�tDA����W��H�[D�ޥ���Q�>����\n8�z�!}���@�#n(�N�N�������\�ך���<���%���3��?m]�QM1bW�����d���xL��vnYs���;�n�:����,�P��TZ�e!��#�;t
��꤭��vf;� �=e+�&N��ߺ��QY�D:��-�p8v|I��N��˭�7i^ݱ>Vf���j���,�E�u��� {�N���pOVb:�2���czhl|��YpE��+�DG�����3��[#����*5�f�'�fl�d��YZ<ȧ�z�͸��q�3k���mg��!��!NC��/��9�����F�>w��Yғ9�={�l��,���Q��Ϛ���wޓҭgDP�����1�����V�1M-0��^�e��/�:�HZ��beQ#�(���ǧ�Π�i���f��垣��	�P{�B���9�('�"O@9qX��7�� �W�,�M� ����g5�I��r��Y������٤x�P�[��
&�h���ә�bU���;���HoHg�į(�W�c�#����`1�{�� �r�̺D#9{��<������"����Z&���r�>	����M<a��}}7xh.C����b[;k���3釮�mԓ��aL҅����ԯ%\������n�9v�F$9�56�n�dY�sq_SCOw�UY��?� ��T>��\����F�����tE�|������a��N}�}i��&3�Oz��AY7A�Ӕ�/���f~�&����2��N-�H;�(��IÙ�!t��Uؓ�{M���hM����e����ʙJ<�m����3;�H��
R�+̇
��??�̵?�ߒ�/��n�:]�9��h�� �O�p�l�V���E��^�]�mʨc#��+1j6p���S�"|G8#jf#�ԄD�R�F��x��d�;�ɭ����v5+�z����Nk���fZ-۶��H�6�O�J����V��[Ja�q��3��e��_�����"� �[�:��|��?D�D�[���=��|��:�0G],�B�t���n��M��v~̮��G`WnHY�i��О'\g?�! )ίR�k |㑶ё�9��<E����?��Or� 0�T~y ���i�Y�R/dy<Z����j�{U`(�W)ǴGv�RW~�ǅ"�Ѣ�*����R�e��n���M���^�Fo\7X����y���KN��Д�Z�
L.�7�a���ڟ4 O��G\
��{��7,�u��	z^S���O��I/�w)[���5�sZR���c�̚�C9ק�ք���ҡI4!��!��D��7�Ɂ����-�2�]䶙��Ə>�~)f���KU����8�[-�ЃY��� ��������$����f�W�8�p���m<_�G�[7�A��P{O.|�~��#��ik�����bʨ��Z��T���N-ՃJ��U���@�CV�-�mP����yU���$���,A�Cl���yd&�'L��=^�Z���ħ�G&.h�	4�ۍ݌{��z��0�f����*գ#	�>��c�sP��
O�s�F�����R�s�����ܡK���b��!��r1�D@�L^ɔ�7k?�#�N-��|܉��]���(ғ42�y�T".�;�"E:���3���܂yŃ�ό�Rۆ��s^�}���3T��
�uG�����_~�p0�n*�ɔ��pl�K�R���`�H �gT�����	@���*E ܇���2��{"s:��~�}V��?6�u�AKW�{@���Xv�7
AivEQ"��B��T������I�I��]'+a	�L#����U3c��Nd�|?Aw*�E_�o��F�A(]7�GY�#��]���U�:�v��.K�d�1�@G�ԥ�9~���H�G����]f�T��r�O�3���O�����%{BU��ղq.�&K	��v3c��\Rw�fH��b�e��Z0v,�l��G cP�K��N���<��:z��
�Fj�!�r�(
��;p�S��D���x����k/��fn��8���5��\��Mv�_e��sF��\SM�r�X���1j�k������*���=�N�,B>�:�5�欏��1��Ep��۠y) [��(�:�O�t X��_z�%;~+
����%�F����y��A__k�cqm#v�c�	C��!�8��}x��ܧ�����%��V����cʲ�y�/�����nGƀ@m&+��ے��7j`���QH~$"�_��UD2m��e(I����"����he/�JC�5ߙ|+��S��L%,Ĳ�	��v���H>H���|I6��|Q�Y�)DTd��ĭ}Y,#~���2�櫣�VXp���U��!%Q�L�\�pa�U�p�#*Ue���sx7���$�C�r8?M��)��X�<�J)]����������\��8ȻBվk� LM�%ߣk��h��Q�i='Q	�b���s����*Wo�R]í�j��܍q�(:�Q�	(���c}��1�*�|�&�A@����T4�i���l�����j>�o��L��|��b�����r��v���� �~}�>��yL��C��SiO"QOӛ����ţ��E`�:��_2�|���k"�+g>W4(-�A��1�%�pM�uן�X
��dC#�ϖ�&�S��0������{���5
���FSE\6pg��Y~ Vxï����Ȭ ��H!��{R�5���]G_����%%7ɯ
���S$�s����/�/ȟXw����P�x����6^R��p�#�g�<��p�fc�]�f3����4x8nW{+ X1�"	��Y-��2]��Pĩ��n�)*�f��@}��;Y"L:��kj0F(�%���Q*��}�Ñt>+L��dw��hB�.�xEH�h��e�D'�CRU$�p:�^I� ʑS�7������%C�@e�LطS3�f�Q-�ρ!��!��#C �o&�R�=������r��5k��^��?H�ȝ)�$0���o� �(���J1���N&��� �`.���H,�~����q
�K�S=��FW6F+�C`T�$t���	!`�0��@�\���$�,���:;D,&;�@,��!h���ޕb0<lO�7�s�����T����zx��{��C��z�I����%䤇1Ek�1��aw�SWm�|�S���Iv?�����
)����7Kα���و���=�
��k�#T����e(iR|_9��P�Ng�.��+:��g/-����u�;�'C���=�[����k�Ơ��S�S�'����[��K�CxB�G�TX�K���³̭�`:�V,���^��*d-Y�yD�s7����l@ �#�m4V���9�{铌�]����j�o����u7�I/��4�q�*5��b���r�k�i��L�����ܔ�WV�l�J��Ƚg�\\�'Hn��Ѫ8-�]�����5^��o������.x�*���0�zof��6�XoQ��U��f������6� [8J���9"v���lCe����A�97Ɲ�и�u���I<=��	�G��O��f��'���)�ٯb�R�SO3;���ެs��KE���oW���v��p�.�J\W��m���h�N�� 9X�71g�d@"��<\+�=(�2�}���~�|#ub+!�i��_t�������K�2�>.pu�C�L�*�w���"b�>�M=�0:��3��3��4HdU�!?x������X�G�oR�zҳ0���5Ĥ�P���#R�q��
9��������#i���l#]�� �NM���
ڦ?#j�>�	��'�= (��*�6����;�D��!�����:U�Q�ZGm���c؜JTm&h`��м1����y�69���&ȜV�a�ʨ�`@�V��{	}wD���6��.1�;W^Z���l���-�����"w p��d��4�3��P�߅e�x'���q��[�
<WAy�5x}�]oVf� �_$W�=^G�"�6C���������<O�| �\�8%������0�|�9 ����	�I��E���+�9(�
� `���i�XB�B��cb�[���HX����<�]�� J�zYr��6^��UX�ށ9�G��j�Ke)���eŊ0VA���&X�
R�I��,X�Ϭ&���iK��o���S��� $!�o�'�͠X~�͎m�����&=��P�2�ۙ̓�ݔ�t������ﭦ���{���a:����N�]�m�Գw��~�������{��i��6}����񛕎��	 ��1Rf��Sgyb*?"��]�k#6�Ɩ���m8��O�b��T�����Y�L��)���~�vu���Y�7��CByO����9420�Ϙ[��ߩ����ռG=���Ϲ��Ph��3Uz�'���̪���`(N����'��:����DJٝ�k0��ju�����RP
u�����Ԛ��|��7=zCJ�c���eOb=	�.����U��������ϡ|�7,�Ss��Ss���#�7���������kL�;B[���2՝�0V�m�\8x��\���J�E�l��i����$0HLCt,��#[�YvE�.�!f�J���]��H���m��D���ٌ�v��&���d6�P��>����Z3%(�2��ܢ���}@�q1@I	�QnW���A���6�4+����d���T[[ycJ2�z�-�W�V�� NU�jL�&Է���l���j+i�#��)Sa��_��m�N���]���7��=6-P0-�@<��a�z��3�݋�D�]t�S^?ye:�/�V�������Vt�d�ݥ�E{�����"�-�ηsqw��t�W����'��D���7�Ή��@u��*߅t�Q}]i:��~��MO�4���'�N�/Ǒ��f�X�[ �i	hmitDO��W6J������|�����<ӟ�����*��xoi�)J��{(��r���L�=�3ĭ��kF'��%d��,�=����vm�7�ꄲ�M�<c�wAS��M��������00�D
Df����o�B��K�¢��Q`�Fsr�m����7��ݞ�We�YAxn��@��{�}�EN\3�ァ�HN�W⚀���z9h�t�k�c÷��\\��<ɫ�O<^ρ[�,yJ�W��*ȫ�CH�M�Ǫ�I�4S�g���hd�?�ق0d�@���Vq�Pn� �%��mlÌL	;�o�����gA�D�2_�Pt�����9Ʋ�B�/�X�Tum���-���fE3����?�4����\T�_����Ŷq;�x����3.I5���.��\�{��".����s̓��-eC�+@E�_�WD�:W�i�c��,��T�W��b��!U�i*>0;�V�5ᖤD��q2��� �Xm�&����Ҥ�3�����ڰ��Ė"h欫P�RfU�)|5���x���`�൉�~�kMk�cx��K7[���̉�'�[���y��J �fٳE/gϧ[����5���m���{�Jͪ�&�{E�h4�	�����Bf��Gz?��[E�Yc3B<��5PY�+��%�'�\4V���0WK��U_,�i����۞��;���h��Vv�]�҉����[�u�W�Wb�A��o��]�qh9�}Sn��<cF��$bof�?�����%�
���~,��i���^�3�:s���v؜C���R���<o��XP�2=J���2=��b��O�#0`�|@�:�7���X�7�q?��Ǭ!�?��ږ����ӵ6��>��d��1D�f�RݪB�
�u�fbl��dD�N�_·}<�P��Δ����=����,�R  fO}#a��\���ҙ�)E0P�>f�#���x�|��R|p���8�R�B��YRZ!��z9��[<�|8��{�9]Lp%F�+k���r��h�nq%ڨմ/�)������8sڵl�p���xe��Y��R��n��h��R��S�[�������}rI�.����&��>Q�0�a9�&�ֈ�/'���)=X�Y5��+��;�J�o������)�Q]6�UƸ�6������=�;tQ�6d�aO���l�)�F�p�f��l���؜�CP��4��f_�J��|$��~q��LG9���>&f�C�����v�H]j��X�2bK�����f��E���x�M����3~�DH4�$�l_������x0�Q9�]Q^bB9cb�L=m�|D��v4���g����9wO�z��32��]�A{~�ҋ����t����+���'��AP{�9W���2�����~}Ƒ�)�&d彰�Б�@:'�c���b�32�>����I��+��H^��Q�9�论K�6^�	���tI4� ₒ&��P�|��.(����B�B���t�˩J��#����l��l����<�l$%�J�vfx��{��Ž���}�7�"ֶ�ろKކh�yWA��M�۟%��Ϫ��UYj�e��|R�$���NC�t�G�Q9���o��~]������X�"N��H��K�<F��;���`�"�����@}���2!"��7[aLec
��2��.�=2����VG�bɍ.Zk�	.�0� V-
����ⴰ��C����"���c%��y���X�>߬D9�=�rL#�%qEF�y����fF�����Uu*=�g�^�Xcɛ�9���5�@��;f�g�ؽ�������T �vc�,��|!m�`4 ��DJAf ��=V��`�u�8d>Sh�qԃP|�(��
��%V�ko��X}OZ�\Y�c�$VBߝ� T���ęl$��a��$FQ�p��<}ҕ�R�o��������g�\]��f n��s�1v�+V[jH��:eܶO5F�b\L-�rEj*�y�t�{#1�����Àu%>쪧�e2i�f�c���+i�[&a�f9#�G]����B����CЩ�BP�R��T�̱g�H�٫c�&I\����6t�����C��Ԁ�f�ú`�������c N�M���.�v����"��f�S���Q$��O����x��>y����g}\.�������@�]�-����2f�pzT�?����#Z��֖Ax�� ���D=��,�n���gUU���9����S���q�F��#M�7q�\�h�(���/p�`d��H(\4�j�&�9�� �U䕭��w�7(���a������?��F��R_-�4�YzJ�^g4�����~���@Ϝ��^��H���)��#B��4�)���d= ��3�3g����
�j�Oл��Ü�m�?�1�9F��/��@���Z�+��T�8����ط��^֬�t���ٖǇF���������u��^�����d�섲��s*,d�2�w䰲�FI�����a9���+ ��Ɋ_N3|�$>o�8}� @+�"j%q5@�;Zf�j<7���D+6I�,H�k
ӧ���@�g�ut~���e�!��t���).Z]�K�
��1"�W�����G�se;j�����t!׵s!�v��HÒ�PC�x;ʰ�ڋ;���?�|��ۀ&�iVF�M)Gz�J���03q�+a��N����x���A���1���j���f6�X�Z0�7ž�Ue�>��,���U�p�o9Ly����A���`��X�t��s��\�&��؎T��9z0�N#ݎ7�Y�73_�jm\�*�
$N�IL911�	kϫ���w�����-��ʶEM?;��<`D�JI�=bO�pKQ�mѽ�f-�3��"D�E�𫃂S�#6w'���21 }�+�kQ�<B�_ZYF�5{s����c�
���V��ROuS��H���!��j�!�3
{q7��'�EU��	ǩ�GF��Iu��Vebz���j�qr�e,�ܾ1����6�@`�d���=�n��Jr�qҭ��;�=�Yh���A^�0­}W�d��n+�B&�#!B��S@����b;ۮ��!����_�	��(��I��LǗ�Zm:Y��;r���eˏ /2N["�l�yͨ)���5[J �v����s�Q�3�G�y,��ki�,>~I��G����ځ�]��o�2fyܾ3���,��+�¡���8�i�%A�\�F۾�2O~�I�����F���<n�N��N���CB�����Z��Q�ҡ4���(��Z��G/�����cQ<�.6�hS;Kɼ����- �5��,H3׮?ɵV��/�g��%ϺA��v��#8��t�D� �`�rz�W�~[刎/��x�$*g'{s&���z�/�i@��A��i�k7�dHa�/�nE�H�4;~�0�Le)�F̷|���i>�ҼQ��Nx�u��C�����̽���=��HƯ�R�A6WhU����iݩ٩`����bˆ��m� �H�Vŋ��z_%�^�tt�Jz��;��Eԛ�j�Tq�8˔�K:ukў�+uV~�nA��S_b����gyC�~P�l���4�Z��h"с~*�����C�>��k�\���n�zO�E#�Ծ)��S�{�f�\����ߪ���ڶl�/��\��/��9�R��x.C��9��F)����%,�s����D<�%u��d�@Yf�Fk�|�E52���I��͖�`?e����l-�0@1YS�*=�<���B�5��A/*��}���Yr������U���q���7n�?�14��� �G�=m�^Q�R��	��Pύ,���;��Cq�];�FSK����S��T���5�-S��u`1h�S��+�C2��{�xQ���U,�D�[O����՝���¾�
��3F�`3Ӣ�����>J5`���|��I뱣�=�^%`��׿j?�v�NN�!n�|3�f�`�%2fA_/c`���Ҵo�	Y���2C$ڰ'���Ñ4���J\ܺ)��{$��m&X�����T�@� �W���S��k958�kR�����%�7��zO�s�*7��E�K�R�l}plLt��5��0\H+b�����0�/Y��vឳZ3a���zP��;��wO��l�m�p4�	��!/8&^i�!	�tdD��3�H�tԽ�.�d-�<�D��C��'o7q�\�DN���T���;��q
�b��]� �>џG_��EiDXE�能�%#B�
�lI�-�:����F���CԶr�{�j��ف�͋qB8[����}��K�Z��_h_م�b�}vLt�eZ��ͤ.��OM4{T�f�\&�:��Ot��vG���#k,�������&(8mr�7�E;��������A�No�"z���$��>��:e(!��5)�潫��i��)�@M��YHe�j���g8L؇�r�ץ�/��?��#�q��L���o�ȵu� 3'� � y^�7�Q)���I����qŁ�Y&�v�� =���%]s���\)�lۛ�K-�����@��:a٨*h�	5"��I����T�� ��eZk��l�p��t�V�
�̅��N+ ����S/�����$�-�;��s��+�]/7�� @ּ���ãPQ�%tp��㥼P��L�8���1�v�~��2�)UH�q��hGH$1���C{
���:b�B��mNT�M�����pJ��@O<t���b����Iug yy�yy���b��cq5#lϣh��rlS���pI�ϯ���N�@0Y����K_!=�m+��a���^�z٬��&I�@B}D�#���K��}!T���=#�l>;�I��0�Qtg)�.��]t�L��.����1&N��#��� �ɣ����2�p�F��}ܑ*�Naw�i���&�2Y����ɨ�9��4���!=���c��|�<�@��5��``�~�8�6�Jz#����x���wG�C�ay�2�06�Szw�쉆��)�zpF���l���e�x�>��Or�.<
NM���[&u$�[��T��΋#�T�Bȁ�0���ސ%Fa�����ϓM�睚|�w��xq�R<�}VrM�[na�����`tݣ��R�)���/)��3�A[��w�r���Q���k�3C����Y���k�{M������4=��^_�ĵ�KR��Xk��k�/;��X�BCVT�O�{��='�my��xY��V�;�Ţ�[���������T!��B����l�δ~BUx��2z�,�j�A>B�7�Ծ��,�Z`�؇H&�c�d��S3�44���Q��q
��K�)%viYOg(<jI)��@q��qI���Ww���4�Ӄ���ZꆧVV��^��c�b�,%��]��|��tm[�W߻�j�
�6���D:ڄ��V8�1�7� f�`YzG�v�N�
Dq5h�����^@�	�Y�C4�Rw
\[���8�	& �wfW��+���'�T�ΦT}��u
A�t�����H��!�� ��P��zp&��(�m0���2�=�+�2�v=m!�]��v<�1|��plL��ͷPb�מD�wס����c��B�0�)UX���T���t6b;��w�P&9:Ϥ�F:s�W"]�j0���~���^\�荛}K�N�|��ȓ�K~����#��k��Lw2������_=Fȓ��y�ƙٯ�����܂T ���JW��8U�2Bj|�A�fnd�P?XD���Q�[������k!�H\*��%��"�{�kgk ���q�ED������f,���*�?���m�s��sუ��W�T.Y5���'Ħ�<3S�}D�毕i��%���g��R�� B7�¡�nE�x��ڄ�-#{�/�ﾾSm��ۅv&6M���NN��ڡ�= ޖ��gp��OP����5.�-�ƕ&?YokI���7)��h��eP]v=���L��To�Ţ?+d�[!��}�U
b����*rg�
�u��>[*���7�c.���L(n0�^�jW{��	�ğ%�H�b@��<s�QD�h���DJ���7�8��+���π���T��)���e
�9�/u~�)k��͸�2H��7�Y��ۮj��~�V�BZ�nC!�`h�u0k
������I0��.���\�%��GX��|��+HJ%]Z)�W*,��lGs��$3�;bOg�a���(*�y�F��_�
�QS�0���T�W��"�&��@��2*$j�áͩŪ��2���l_4��y�ge)������S��#p�y�82@�}:����_���'��ֽӓXi>\��1�h��_E4�7jRi߼UH�N|q|wJ���F�����&�(��[ME3��;|#|k���%�P��
����&��	7���o伻)�*ۃC ø�E���*�z����:��ǜ6ӿW1A	i�3*@���k�:h�eӲ���|��]݊����&�/{{�5�r�m?(�)
J]�x��8����k ��ۥ�ъ�Ch��w���B���D��Lz��ط��n=���{���$ 2����X+ߚh���@���Yc�Z&���^�t"pH���&@��	J<�5�L*��Y<�@�C�0�V�ԥ�>�d9��|utu�I0�@Yo	y���~�@��&A��}�,U�����Vo�Hc��˿#Q6�(X�ǀ?�w5�%��?�7���x�WC'`��)co�r������[K(˹��?9�0N���� �'�c+M��r}�@����ڼ��LoT��PW��Bb墵���&o"N�qb���\����ڹOBs��%g*���,�"�1š&;[�ѯ�-�	�8��[��g�pp�Ԃ��K;���
l��Ö��ݢc�B�Va}�	�HѨ��PtE��ʛ��1}��K�De«8']�:3��d�D/��ӣ����U7 �E>㻤B��L#Q\��x.��0�~�a}���S�V�K!�̢�E �3�́a#ޘ�55���C�OT��~��rT�B����eJi���J��u:�%��Qh,Q�y��(K�8�]��Jl�r� 4���^�0�ɢ1���=���6%_]�-[0�vb��#6�䑥���T$�8ر��y��{��S�~z������j`�N�'�����%Ӽ���@�)�x��̾݀u�����WH��ל��T仿�dȿ�4�	L�����Cmǜ��V;��4P/08��R4����SA�AN��
���(��u��P5�r1�r�6q�������j��?d�[��e�^
�AC��J���\ȧ��XK�����v�i��p%�K��U���:0�8��q�� �g���]�!D���c�O����ge�Xk�V}�O���rd$ڪ6��J>��j�BJB�]�ht=�/R�o���,@���I<FpN�!��R���<*3�2#�"	'�K�me2%4/�2]� �'���]c?8�)�rH��f���;Z��9K���LOt�LЙ�#<�f�Z�U	���Y.�})��KC���`��%��W�����_��0��'�x�s�1�:oQ7�<�oe�Y�{�����k�{�V��q��w-<
��d�u�������E)���6,$�zNې�w7xP B�}���'��H���b�S�.�$���< �^ae~
�=v�[Gv�B�	�d�M7!'�R�Z�!�<^N���wt?T	��?�b�z�	%��=Nba��~��nzx�4g�T�z�(o� �v����
���|�U�6�GV��w_�ՠ��PB�?]*G�E���/������8'�#�r�`^KN���/�F6��Ǿ��� �boެi=�?�5y"�!����3QR��w�M; ŝ������s�6��#�T�C�N��1�Bq����>ƒkr�dت��^z�q<��:����^˛��Dp��X	�M�E,�I1��8� �E�P��EO~h4��jk��Q7�%�X0MP�-�3V	�?D���0�;B�8��Q�ͧ`��7��K��+��s�wrޢje���e��-�������SC�����m"�{㎝hu�s8p�5������w���������
��Z�^�V��O :�����+Ċ/��9t��� ���<R*ֺ�*����;ge�69PI��t�l��2V���jPP�M93�Pcx����N�+�� >���>=S_�7�㪃����؂��V����/t�����	�A�ٴ��?��kɞ�Q S��꾻SL���x��o�!Q�CvS_看�:�D�f�:�<i�p�0�V/�	���ҁv�B�pMRV��wz�T���E53�(�s�ryF ٪<�ğ"�"�f�F:L�o'��Щm�lye�7`=e�d��1��b�!̑!|�!ށ�v֘C�c�����`�#��u�D�V·"���+�����p��aU��xm=��k�~��&SMGT���G�T`�p�AӖFP.>dp�y��kT�d�:��\���Bߐ����B�cg���>�� Aa�<J�d�'DLщ�~v�����k7�����c_��Ua���D�:L'�-��Wm�P7Iz�W�RY��/ԕ�gd��A�� ���tW�����h?[GMf��/\3��m�����q�2�o`�uRZ��W5	����1��1��*��ف���I�hiYv�W�L.�%�5@�o��O�z4lkܦִB��c���-��b��bl�]��1���9��r˽]�E��D��
�½gP���o�cHC-	�OՏ��� �%�3S%���:Zf�Q#�}x|������ T��/�,��f)�pBRv�L��E�vo�x�Ok/�?aӐ*�����/���b]C�6rO�#�ۨ�r���W��#��K)Q����~���ɳ�Q�|���#u�c?&�J��+j���0�P�����G
ױ�MŨ��w�Q��W��f�������3��+��G��HT �#:lbGt#�JH��nv��`�O���gp��L ̈V�g@�3
��7�IQN�4f,n�}&;Z$Y���I�4�;��M$�.6����R�~���i 
I��+t�+r6�6|�T�������W�4}��uq$�5�`��K�`��a���EO6|�
��*�¶�a�8	4. �w,x�\�8�"z�&.>*p!j�����&���'N=Y������U�T��º�c�I�q��Ĉ5�|�H��
��@�X�=�ҁ��J��ĝ���e��=�U�S��?G���L���]�T62�?�_�gg�<�	����DuP���
�]-/B"L��T�W�;$�qt���\�x�U��'�t-4
�Q���i�[N`�2'�l'�j d)�ߨb���8{�~�y��=&=�|֒A\�K�rWdhk��e�'���.Ɂ��n��K�]����<��%L+D4�UR@�H<��}LL7<��u\���UϷ���[�iYE=�a�)d�ٟ���-ϲ\zM�ꜟQ�[��r�i�W
VC����ME"GQ�e[���ǑĎ����z��{\�[o�JMB��6�B��j�NL�.��;�����c����������`M��[��Kg ���-Zd*�����%V3�����r�b� ��*&�v�����k,I��@����c�?�6��r��yF� T��0o�J��t���ѨXH���P^?J�AwhB����'�~�?�\I`9���SviKC)�P��`�=/��J)�Q
���]��	n�'*C	y2O9��� ��>{���7��+��"ӡ��%�|(i� 6Q�����r?��8���3��ᓲ2P!�(�طC�IW�[tZjԾ8|��<�k4b#3�E!mL��`s?*߱NZ����ͧv�Pﲡ��p�������v'9G
��%���ԓ{e"�<���������v��r�\�r��ty_�d�����p��~"�Y��8��l �����f�Ϳ[�P��D�q̒L ه�!�ܧ ��
CF�Ӈ�+��S����+ ��z�5f�1;7c%�nE8/�S���x�g#�>���<�['p�Jw����Ib�WU>�@�΃rh^�d�q3��Y�D|Su�m/�w��B����4�Gߗ��)�c��l��Ѕ��d��:1���rT��[��1$S.�Q��&s�*�Z�q�1�~���-���=�N�d9&_Nm�Y��@%EW�zӄQ��^$�,Pؽk�Xy�������5*�AM���%g��}�;�h0U��?��uV"�:�*&m�/E\Ȑ�[w�޹���&ZuhY��0$�w܃�t�Ȝ�N�Z�\u���D)_z{�K�_�
}����
S]��*�y��>�*3�ԥZy�ե�r�3��*���M>�A�g&_�m�p6?�_j��`֡%/�c]�-r!�=�/�,�:B�mh�ru��-�%#h�S��I0]�&���ꐋ�אh��.� C3z-4�L��n�^`��I��ų��g�̋�{��ʿ�r_�}�4�u���<q[���n\�9��r�F9`g�u���'�w=4P�3\���Vي�C7�L���(�@������|u<�p �;YP?>As�����"H�V~[�����K��4.�I:�600�(�+qL]A6X_�%���hҳ�V�=�0���a�x�N�ᢧ��:�H(�#[���ۥ�Y�M6�UJ�[����:�,���#I݀kV7�ΟT������(Q�]1�t�	G�SxH}�� ؀�n���P�V��J�}1���)L�9w��kg}�iY����X6���&9��t��� ��Ic.�k?3P*q0��R�fiP6
�v��'%/�Ѵz��%_V��{p��|iI�
�]�?�C��?�yx��KX�b�9��o���]?U7����w\��V�o/�����I�d&��h�q%��cs@����M��|�1´�ة����ڨ$����xC��q!��w8��0�A�������E���x��,�w�������a�V����"!�N��i��xJ�r���>k�D�:`
�j�)��=J���oĘ��{3�\]΄�)e֖EY����P{��V�HQ8���\!z#`#��o�կ��𥉉$��P՝:qo9G���V�']��'|����O�@�)ț5���La�� Z!;g+��I�o%#>aԜfxӅ��e޼J�sQ>�9DP^P
wc]��xݢ�I��qd�Ի8HX�p
8O��6=��A�ˬ�e��?�CI;sR���
�J-��D��Sit�-'�iM���a���T�l,�;�.I��
]�T�Zw�n��E���UfƗ��yU@:��AC&hL�!bj-�]�s	�
{�I~�fs��	Z���SK����l��Dwx� aA��ny������p��]����*�n0\�Kߞ�%�i��F��՞������!)�+1xz����N
�o����X�����Mx(٣���Ѿ�б�U�=_�a�V�q� )P�}����6��[Ǭ���l֟e,�5��w����_nH��f/�;�qeNjލ�3�c�Z� ���	�s�K��
�?>��q��AX#ޜ(���J��l�rX�82;~��%�{R'ґV�\>k|����A\]5G��F@�;|�oh��}yB�Y}s��M��^ߝ�Ъ��	��[7�P  ��M�vq��_R����Y@bD�Y�/g����m�a�B��.�N���G��`����4����D�n��M�����\e̚)�?us�Oֵ'����̢��I��ON	�����S���d������Ä$�V�=Z��@Sm��bM*�r^. ��N)༢d�\Ud9t]wK*�BB�+�l�l���{^��S��Ί�c$��H���8�v܀5t��7ltHߥ����2>��̽��d��V��Q���ʣ%<����8�ln� ��sh���4eL�i����Q^����c�%>E�lV��r���ê�B�qP%�4��Me�rā��6��?44�>��z�jYy�����0�q��gE��b��!��������z��Q���Cmty�+��Ԯrg������M�J%��X��:>:�A����a��W��>���A�w���v�psg�sϵq%˸y^�q;
����V2R~�U#@;�^F�Na"/7��<�ք��p3�2E�t�0������ r�#?f�l�Ld�%��SY=؟���`��Yf�!m\@<}_IROBcC�\�^��>�9ELI�0(;\�\����m���fwzFQ�O9��b	b�yK���j)6&��ՏK'Y ��:��m�����?dV&0/<h��5E瓚�GY'�Ds� ~��cM���>�U?_oL�?Ɯk�����^�7>~\�L���am=+�S���.覈¬B2��S���U'�\PQ��ş>h������v�P��#�%�f���uc�[wY����~]��lಓ.����`�P�eN��$�G��(yr��0�3�ۜop�[�A`	�@���70�C��cj�t�/����	�����m��u��६)ͥҸ���U�𚠚�z�̌z%؛b�Ŭ"۠k٬υ�??�I(R�
���[	�k��sF��B���+�q�$��ܠ���8 ���Lo5��q#G��� �P�PWmv�V��S�;��� 0<=I��vI~Q�@�K�]>Q����Q�N����)yRppV��P���2�C7Ư�m^J��0�d7)̭��H�$kB������	�����4I�O�ҿ���K���:�I�@�4�	�~�\t��^w�8��̟�(�^��$�^���_ �:��+�V#�F�H.�֡�W�Zdf�+hc�nA;ĂO׬T��O�Pn;�(�؃�����O�YSO��=�4��.��v���	��c!��f4�H�ٔ�����J22f���;��� #� ]y��3N���k�gQU|�qf�*t���t��g:�-���������y"�2�9�bpG�|��"4���#���f�et�ӄt�-P|�A�n�:��o!<�d��+��Ȋ% 62�N�I��].;׵N@��+�:�����;�{}�Kx
�fkFBR׎�w���|��u�+��0��e,�ʳ��>sNb��;�M�6��2�jGD}ˈ�qs�6��[A/ٴ;�z�(��x���s�:�+����C|$p'��;����_:��t���t�_�b�h/�Ta�"�M�BgsՔ��=���]:&��.������r����ZyTT,�2�Q�|Z�_Ef̔�{����#U��}��B�r���L�1X��(���1�0�=<c�Ώ9�nJ�o�߹^^�8~}�1Uu���Ǝ���8o���p�h��ݓ3`�m���eߚ� �Y��ϜX� e�EK�Ĩ�m�q�&�-�T�7�IyG��1���i�]"��{_�%�I6�!���#�����o2�X��>ÕC��a��)l��fn�4 X���W���W�yT��~�RN����+�����
i��J�)�K��.��`ō�9�V1��MD
<�X	��v�-���$�����G�]�������LOq�L����,�
n���/V;�A�Yz�܅\����N��p��Gm�n�Eȶ��ax��yH�%��f;4�5P��.��u���=P�I�f��X��D��� ��<�xwX3�[��ps�:-�K8w�%�D���L}^�����#t�8I�}E������-u�D��B�y��CrM�[�j�;�3- |b��JRȯo���;s�T�za�l��t]�釕
�^�YH�ȟ`qU��?�t��3�А����2�r��EG����\#4���^	�ѯS���3��0c�1+��ʃ⟖����QBl\�+s���v�kl��W�2�$�1R����}�֫�2$�xd��*��}�;>�_H'��h�{���!Rw�JFG�ؑ��Fڞ�¸�A����4C��@��:�m��T"+0K-Y@-�!<�&~d��,5���Xy1^��O��ŀ|�Tg��B�m�c;LBp�͘�MR���\�-�|���$�Q碑(����G3�;�n��l��)��������k�s�d#4.\���n:Gy��g|��e[���������������QK��(7"�#���G�E�-��K�����S+���m;T��L�����<V.F��){����K��k�`ι16����v�h v���&����m�RM]����N�:סc#�%���!f� �A����T�p�S�5��SVg�y�`�^����5�d���-�:L��!�5�V�V�~*i�/��鋅]�9S�����tm#�`p�ǲJ�f�����タ��)>�l7��� �eo�Iz!N3�΍�#D	��ـ�H$ԨO�/��e�1`���X�
��7�4�Ea%@��v��2��G�<JE�T�J�2��~Hw����5q�� -~�>25�d��Ku��ʆ6,x�/�lI[}j�%a`��IsQ%�t��k��r��0/�,���)֏ٶx�+��=N�s�L�.� �[�rL�з�:~4��gxߡ�(��T�	��w�?Rř���](��!�\W��bp3Qq�c�>�3�Zg_��8�S�l�5W������������Y׮A����4,20F�a�'E�r;p�?�'Fg�D���-�y��L�1Ǵ0E\��.^���d[)�̎���[�N���H�t�wx7 ��Dp��E����W���>#w�{~���#,�%�Ӟ�L���Π��5���������6�%��Q�B���5O���Qxs჉�~-Bv�K$����L:�;��Jxn����Q$�����}����#����M�UP���hM��[/���9:�WU�0m�c�n'jf\/:c�b,FB�.1���
$�ҡ�0)�Ǽ(�5�o��'QP�a/��tA�搄\I�	��/�:�ƪ���^̻�y�MR��N��+ͤ_��$f�/+��������5]do��� �'LF�l�	w#.��#���YV"���m6�1D�qff��8�a'j���h��À\|]E�z���E�g�"O��,b�������(�y#TV����y���8�+���?9���SyCŌ&��B�O&�_��^	֘�="���M`�w�O�@3�|0:	�ˑV��w>؋��^5��R><��.��"�\��5
�W�1����o7�DfLv/� Ԝ]J��˵��n��w����j�8�ރ�t�$���k����
�6��c�����[E@@%F�v���g�!�4�(B��Ӫ�&W�\��C]Ǵ�{��#�?��E��B(v�ne��� ,�h���ZH�� i*{�O���2Ш����k��KKWe�'�΋�w![rJ��7f����%�(&��m7�ΐ�w��5D~\ԐɿEĹ�ҫ�~%�t�"���w�U(K�̒�N&�KD��� ��)��kB-�@�t@�]Q�O�&4���)�y�:"fVw*Vcכ��Ӧ�D��֚}h�]�u�X��oV������.��(���k��Z����1!cq�a��Y�e$��L�����+�	dG�
h~F�ag�
�8������r6a��� ە�J�G�/I�	��nmִ����e�U��ܚʙ����{��ܝ��z�W�M�NA��74��D�V� ?;�S����6d��'O%���gm,N�V�
�{��/Q���z��������F���}������l��~Y`m�u�T��`Bv�V@���K�������rof�8@n�J��^��GE=A��?�_7�e�]�&�Y���:IϧĒF��Q�ڳW�`�� �B���H��K�5K��g��x�ж��;1��wׅ�jU�$fB������Ækp�ZB����I��(����⒖08A�ش�J�7�����_�YE��2jΛt��bQO��/��`����L�{�&�U�u&��ZS�~ ��L�et�7+;wϵ�m��k�hz=�j��\����a��.#�Mm��G��i/�9#����~��;�����n�Q����@���!��� ��MIO��v7���8��@��U]>�H��'2�H�-��e&`�L��w��6���K��r�w�ѣ�j��Q�Y�b^�5�&�)����=� �6�Ek�+Ig}z*�0�*:6{@�묑" ��!8u���5Q�a�����>�I�Ȉ9�I�g��\�)��ϯ[ݿ)CĪmJ�O@]h��\
����	UycH|���yoG�T�,$p#y���N�jħt��g��5#��{R)�ߋ��l�	Ӝ:p�N?�MY�s�����<�ւ��"�e%���6��]
���R~�ӈݗ[̱��v{U��b.�&�9���FOoBG���=�wt�[m~ �%1X��:�^ra�GJ�O��C���Кl�F��>�r_�H���g,��`���G�g_>dX�s�:^�f��R��p܃Ƥ`�?K��ԿC��7�K\2��o&��4�1���
�y�֬��W&f(��)�Ô�/H��}��:���C�	�`L�[�1<-��rr�8�v�J*��_^�/�O�l?Q��2:u���3��5FM�3�H�� ��`]tM{�:�>P��%-!�t���"�����Æ����E���� �J�D|�JwT�U�2P�%���W�Gh�F<_�N�8?[�g��)tM�ˈ�ϩ]��M~�t�ga��p�
�i(_�x�z-l�\�J�[n5�J�Y!�HVb�㮶{�q���FK#GU3�_�?�'&��K!�@����&��yC��=�� �賷�E�*cv/O�V�_��^�� `�0<����p0��u�����J����T"�=l�v�L2�3��b7�`�H�7�g>D��\ \K��?�N��ht`��[=�I��݋��p`h3H>���dWkr~���!ڤӲ�^8C�0�R;%X��:���&gJ�6�ey��oV) �	?�� �-Z
Q���k^�,KΑ����h�Y���K�V&I�A
:�"-�Iɋ�[0����]��_+�'��S��M�B5�4�(d��������z8ќ�%��z��%��N��)�"OB�g��]&3`�I��zn��8;ަ�H�1�}�j�h N�s�Ñ��A��	]�O�vQ	��
�Y��ȿ���;L��Ӣ����ma�6�j�(�׷�=p#��,������$/^kl��B��'�4��p�u�^�"�j^l�1���5������զ|�)��خӎ����l�'�t�w�q�nǂ�p�(-���\i��X��Yj0�o�Ǫ�{bQi���C���,��r�?Њp��X#�x�9T�o�9-��|��5�Ѐc_�E�w��F'���\<Z����`"�-ܥ�	�h�b�c�\`+C��V�.�xz�k���B�|�2#�Y{E�#jA���5�����m�\cU�*��3>��Mݞ��3�o^區��&�D���zB�ۓ���t<?��keUF�h>��A�=v�H��P�"���~���id�c�	�sxͯ֋�	�v#h��n��h�# 6�g�.�t8��D��׷�iw#�w�`��K�2�E^|˻tZ̑�kyh�����U�ũ�邑�V}M�"�s�wtv|�����y���L:}�8Bf�Ӷbb:G(�d���(U��Ěs3�S�Vs�c]�Pr�FY����(׆)���_7�m����hd��@	�ĂZ$��xԭ�b湄��s�,��/_fǺ�(},��ٵ�6,�P~[K�����ڹ���Xj���f������_��V�7����,!D�͸<�RLVR�٬����~5ww��uD*�ݫ�����D`6�ӕ@=�zc�8I��@׊�+t]���%C:rжӨP ��7����G�z�Pr_-��!T\���O�˘�-�h,��#�=�|�g(Kel�C:��OT�Cy+��h����j%Ki@�=t�~	����~��W�D{rR�͵ZX�����:��ue��hҶ���"}��T�����v�I��`� W�R^TZ#�9=��`����!�}q�e���]NS�V�)������ҎO
f.=��`s�YI>�Sh��)��(+V���7UGs>j#J?]�g��孤=�ne�����	'͖}EZ��a\�Buy�I~��/��78%m8�Y����c�h��c�;�0�qr����͹�l��XC�cQi� ,� ����e��6�aK�h<�.ΑW���Ϳ�9�A�pM$� ��I6��j<}C� �3�?����<�x+�\Ef��<_p�U;�K��u.��v����کؐ�s{���r���<#����xsAȮ��@d~�
������6I�w�v6K��@MX�gfF
������?:���E8���.r��Nѹ�O����n.�+�33�Կ/��e���p����p�7~m	�=���a�FTr��rg?T	��w���6h��*�J|o���Z�m2�/��M�q�d�h�N�~^�.�O���D��]�D@��J?�Y��%U���/�8mcu����mlT�p�7T�([tM���4�l�6�W1�ZwS%��`����G�9��s����ԉ��M�������Dr�XB��(uU�ʋ�s��#�m������9Je�=#SjzT/9��G������qз�*>[k:���3�8�L4hJ��+�ҁ<r���gP��W�9L��C�%��q6��l�k����0��t�Nsu���5�ջD.T����x�ǿy�rq����+��7np��O�I^]�K��f�	�Tl�q��ߎy���޸���*v~�q����ɀS����S�PS�����Q��EIVs�� ��b�S�4B�n�k0�F��D��n�	������~���Ѧi͇qP�e��!���%�����[�!5��� ;�;,ߺj� i�!��_,Q+[�a��+�¡�~��TU����΅��{��YT�gd.��G��ޏʅj����N���eb#�#!\��qA�V�8�X�>Ԑ+�^D珳j5?O(�F���Y��s�~�Oh��sO˄)㔌^6^�����1V��=���K6��R8���i���V��4�b�7�INk�f�*-��
���W���.�N.�G��lX��{���A�7��;��=��,S���^fv�3��[�&����zφJ��Y�ZE� �,������U&z"��<cYſ6�u����ù���V�(ui�8��y��Iz&�q��G,����F�iu��N�G���f��"�>Mt�>��N���#A�r8��HF��
���8�V���։�������BO=CP�L�G���v�E����4�E�}@���᛾��)ڊ�n��T���*���	��0?G�.>˗:�G���F\{΁O\2挛Z�8�J�;�"~X�¬�(�UIF��U�V�ԁ���yo�:���	��2Z���K�����?��Sn�3�Nc�Ǡ��n)G� Gw��je)�l4DL�Y�	��L�Ҕ�׫3K��V�J�߾T���kyq�Ad��Ј��X�e2K�L��Q�ǜ�S�JI<�4�
��xM����t��{��߶�̦��?���礏��YX�K������	��Sĩ(���4��i6��cv��>�zR(Y4��:iU
t(x�:�oh�.��O|�� ��R"8�S[��9j����N��b�I��y�����6c�遏6b���)������k|O�H�Q�~�X{���
�ib5�3��m�Q�m��e���ߥi�%v�5Iv�k�`>�ş�Щc����*M���ւ5V�+��CJ��^c���
!*u0U#lӮЅ2R��g�?n�4�c��I�s�ٲ�Kza}1D�B��n�����4�^m��Lv `<Sr|j�:ē�ih�VZ׻o�v�/81f���E�J Y�C���u���A
�Q57Ct��᲋�8g@:C�F+">��G���ɕu]	��q'�Z��.��Z��%?�ܩ�ixJ;�iѻf�UD=L��(���{
��(Z�?�R�7�n�@[��n}�~=$���*,�e�K��U�4h]~��K\l�1]L
0|�֍�V5�v[�G�5��3m�g�0��Q�Z����-�(��MH�x�\OKt�b�l�܍Y��Fh�
�i�3S��N�N˕���䍿	!|f��>+	�;;������`�����]r.��Q��1��X�I~8��ܥR�G�(���4Ze������'u�SY���
���;ɏ`|²�oO��/���f�}����x]�laH[{����W�����M��U�$1@J�.[%k��J��_�Z��������$��v����ۏ1�C{� �L��5��QA1��'
p�6G2G.� �9tf���@3ɍOEdlUe�SbJ����Ex@0e��i�Qn\���+s����?��uu�c�	Tvjj�;���9��e{>U����`�a��^f�4rq��69��i���M�ݞG��bu�g��W�DJ��3ڮ�!N��1���f��Oޖ&�٢@Qj�E6�?��
,-�d�w|�SO,%��F�!���TI��*[�֏�ZcHNC��5r���4��	�iŗ��-���q��?7���ޘ�}����s:����N\��[�:�Q?NG2?.z�b�T�8&c��qyɼ��d� ����߈�!ê
�Kɪ���>��!~�����>�!|����%�[�;�k�fJ����x�[�\�����J��mx��w����$]\�J�[{��X���ݧ%sL�T�����۪�.�6ʚ�	�/��s8��;ek�h��%�}
�Ǚ�ݨ3}*4�� ��ku��j;4PS%��
S����X����5�Law��L��z�P�+�s����yӬ�]�&�p�������ӆ�!�^����H��,�G,��-D+�<�
n����D�m���d��VU����}gj<i��P��j��&���&w�] �P��&����v�0��oZܗ�D��_fF���0X��+�6�ʢ8ڳ���H��J�\���$0�9���j���i�h��H��<�Y�;CV�����ϯm��W��ɼ�DT�3}��~M%y����о]S9�����TzbI<��;�AF����-�OP��/�|�
5x!4��k���v�V��y]N�#Y��.��R.1n�#/&�SH�Ky!k�uMtk��*���;~�f�p��]�1�֯3�MX=��=��'����p����D�@��5��V
�p������1���v�'�-Y�N�L |�45�-A��Re�|�nkd ��"o+�;�s"j�Օ�l��ثF�s�+�a��m)k�T����VΩ3����'��s���!��k�伶O1��A���ww_x(�n�F�i& �5`0����?в�[�s���i1���@���$KՉ\�.��G�&L��^�-��w�3�j�����I7MF�����=�~�ض����L�*��|Rmdö�M+�lj-L#�'U�+_��HB�*�Ғ�A��M2$�>/��H�1�(��J��8 C�g�ľ��I�L�:�}b/˺�nP�r)t���kJ(r�`���m�˚R=K��Ͽf��$hh՘V��� ���N�� :���ȱdR��W5�w�n�� 5ڨR��[LCt���i�فkZ������V)N)��g�s7�󛉪��6r�U����)�7W���bA�9�AAA�7������%�=aV��2�,IW���:�8S�|�uk�݇�a	g�N�;E�iF�V:�R�D2�Nŕ�?<�Ƞ���@r�U�A��ܔ`�-��+Ƥ�&���kh�M|4�P�y-�f���e'�a�/G�<!^փ�A�+)��Ȍ��#���ha�ѷ|>.|"Α�0r�	-��
=^��G�
O �t�Mx��(+ul$���Ā�`�Cd��,Ux�f�ЍL��؛�7U_e��W�
�<KñX��v��K��C�5��p�W��Z�fT���*Z����*��g?T{����1�^pg��m�^��_r!+Ɂ�:�������e�nv:j��ڦ���"-���R;���4��7� �gx���n�<�}և��q�1R���+���<}O��ow�چ��p)�;ҟ���9�����;������#�m��E�魂M�¢WTOC#Dp��z{0썝�����7{��:���+�?�QU�Xb=͏���0�E`n�D�ٙJ*t�#�Fͽ��]L��9i=x�Idg@�[�����\Xw�P����jG�kdp��i�q�:���2$�O`:���%[ .!A�����r$rĔ[K�|�tv�4�54���p���l����00��pɩ��!�Źt�I�xa�&�����ғ�H#*F`@kA�3�2@�X�5]����7p;Z��#�boq��t�rO:�p��K𒸚��4(��Y����'�J�"QB�6V�e	�5�nT_��~7w,y��ƫ>r$}�����[��Ǩ�>�ϴ�XʸdK1g�~��e��g;��;r|��C@^Ǡ�F؃��N�ؘH<�R3N�)�3����pY�K \�n.q��?M�P���Z���S5jC�BQd��*:؈U"�.If�[A��҅L6�t����/>�t�����L7�,�N�`��|O�%��xI"_��'ƅ[�fP�"�]� ��E��)G?���(�/OnL�^�P��3P��h��|�a���S��.�����t8�\�ꐞ���V��գ�M�`��:��[aO�
c��ߡ��zs�{/�;_�s\u&�V�c�H]�L�e3N'yҊ�"��أP6頜(Ed�K��6���f�(/s��{R��/�Ƥ�r��ϭH w7�ⱕ�Ѿug^C�fh��f�_�L�vWJ�hA�k3@i��"��Ӭ�Ƞ=y��<�;L�
��r��|�c� `N�[���z|ޖQ?�9L���j���1]�a~�<�O�N":f�Jқ{��,u�,[pcl��-���dD7��y�B=�'RRa����?�:�X�7ĕ������������)"����N����!�&!-!���c�t���V�b�0<=��0�,�|��w�A��m�9D�],��#���x�
/���QF�2�PeF���,$"�B���q'Ƚ�]:��ċ�(��<3��A(�#R�yC��2�'Z���J����*�)xt���xPz|��{8(�zc�PT8"FS������4}u|��g��g�^�_(X�J�@�ãr^%Ъo2PON;8�ߧQY���� �;�:���ߟť�$D��7#i銔@��v>`םgz��Mq��[_�3z�Y�y	�R��@<B2B ��ƸX ���U�h�3s���J�~��E��cd|]ם�589��Ia���}M&r��T�^^\�D��\�2��A`����(_�fvb(�he��ɗ�E^b��,e��j."�0�ɞK|+�����W����s��f�zv.[�}m�s~��oqq�M\�=.9[x�6����˪�-�Y�� i4Ww���ǖp	AӐ����z��N���t�0$ LL���DU�@�t��x��Uȳ�"4$��[�_��� ��)��"��c�c�&���`���>��Vܔ�
'
�K<�"�'�:]���P�ǌ'Z�gH5R���<b)ƀ�5zʵvii2ɦF����5�J�h�'E`݋�G�u���<�)�
��E�(^ދ���7��J�'����5�^p1t(�X8��W�?��"�<�&�
��T:�=/��43(:եƦc��-|���,a���QV��_�yfR��)��SW]خ�9�m2h�F���l��u��x�,��|��&�`_�Ȅ����s��y_˟3�1A��O���nT���JH�:8zߦZ�@�V�m0��&|�`iI��[V���%*K6���F�Fb���Tm�;
mw�9����+C����Х�	j�ҥ�q�U��`��?�Y<u
1b��hj@I,�~_WY����6�h'�} J��]�<�XO�Ó靱R��ۭ��O��s!��B�/����1+��� >�X�x1����pd )V[#����h*^V_�6��as�Ʒ�$����ɮ9���D*'�ͭl�Dmƙ.��ɨ%u�-cR�3�'��&}��n�&��x�>���=���̘d��Z���6�M�y)�˦��X+�Uzd2�4\Z]�	f��b�_d�%
f��$׼��?��TZ��:��/��2tL���]�FPQ{�N�R�ʼ��'��/:<��`�d*���ߤ�R8��͑d��B��U���[US�n7�}!D|����mE�gy\,�TS�k��H���لs����ɲA��s�_�^���nX'�q\�o��RI1���J�!hX+KkA(��R�ѰXD�xo;�W��5c��l�`�v��7�V����,�sJؼdi�ό�ؕ�(Ȯ�K; }�rI�Lf���h�Ƥ��0dhw�� ,%Yj��7A,����ڊ�[;�#��e!������E�Y$�u(آY�E��u�1 Z$��j�7�mZ�)�p�K��1��>����,�5�Dҽ�����ʳo@�aM�T$Ư]�����臷�� �����I�T�=H�����qV��OL�]��M�p�� /L���LW�� d�^�_%@��C=w\ xȪ�gs��R��#U�<�'3��d�:㈦)���L���K��U%h��8����DS:}�=�AG�\\��E�K������\PH���4��>(�eъ��ĳ�qW
�5�u�p+�Ǧ��7I��M�����N���N=�cae��"H���:�a�^����X���Ҕ�L���	������S��հ�p�x}���]�݂~�~���?�g�όJ���oֽ{�����9��� }W������� m?@:o.�������I�3�>���6nѣJ)���/k�^���ݪ^�"�Kg�[`�"����C�o�fFM7NlN�K�����$W#^���}d���nA�&	�������R+,�%�r��i�N��lɯ;�~��C|�a6��焣M����yl�(�_J�
3niIa/|�����\�.�n������s�+yN@��#����%E���� �G�K��LW|��:��
'00-���s��Dج�q��Zn��[�dbb���L!FҪ�W�FYQ�k�[����- �~����6+�z������~�D����e������ɢ���R�*�"�r��f����|�Sp����U�H냁��*؋[��� d^����y9�faW��/ㄟ
B"���P��J�Ҡ:� &��Xqi^�D��Db(����Y��Ay?v�C)�ݑ�?Ħ�M�w10�<}��;����cc�H�(֥�sO�w��&/a"7:E�?����A����m̻~�)X�:�s�w&�����<��
�����>�b����r��Z�s ��sم��>���%��ns�?��}P�}rZaR ��i�:�6<|�]Q~,tC��lbc5�̩Ak�8�1�z�!>��������S+ߥ'�VM�qC���<�<R�F!�o)�xG� �����u�����V�n0Q� h���J�@��Vۗ�֘��Dp�f
��t��Q��
�ox2�i���J/��J��{�o�^W))J��G1 �WlJ��N��vf�>�h6(����w6m�Q~TK�d�[�t}B������s���
B�ȚPAA�~�VdW��M��,}NȜ��J��Fݟz�AFh�^�(z_hl�����?Fi��a�a�5���Z̿MѥQŐ�
�}�~{j�m�������BJ����[x|SG]�r.�+�RD�
K��)|t���6�m�9<��J�� 
�]��΀�=��5�b P�����Ŏ�:\& ����/��N�?肃�XUQ��#����+��5����2|���b����CY��� ��B�S,��Q�;K����׽�;,�|଒�C���N9�ʟϥa�Vr,O�+�{�a��h��P�
<�g��|��/s陁��x��^"0���C�d"�@��ފ4�������ȇ\j�]Ӛ�}�1�Ѷ��%`	J�9��.\�H�n�����&V �ܟ5ٕ�N��',�ie�/�9��=���fr�o�0��O[��cnc�]����}�`��۲��ׯ�	�ӄݡ_�΅2�_�P^}�-n<K���R��l��鴧կ�fOGѼ��e%�n�:w�{IP����|�>�,l�_�%o�+�.6��kn���z�����܅��M� "9mz��7��AW��c`��F.9T��o�̩�X���ᜌ@Ȑ���s�8����s+e*��h� �<�oƍ)/�,������\�렡����bjI@w9=o۝{&��I=�
�M�b�ga��?��i;�HѨ�Ze��C�}Ad�a���冹�3��rL�K5i#�p�����Zw��Co�ccwW�:�Q���Ҷdܫ�o��J�zL���j�W�1�a"����M�o3VY�<I!����V+����햮_pI��T�G�F�9��� ���@3#��BQ�c�h?�ψJ�W�0��TDf��Go��6|D�j,_�t�Ϝ1�����	�=���g32�A���BMz=s��s��@�v�C:��I0���qQ�V�F��-rTf9�y6ZK�2ǫ|��jL �//�7\T��t����Ϡ���8}�:�R �?�*��["®�~��X(��� K5mޅ�B�AD.�,��9փ�J���g���pf�"�ȫW����[߲2�*��>��d��&���[�A��?����)L&�v�Z"��4z?+mzgE���/��:0���}?�A�����L��\�Q؂#	���Om+�&�x�sT����LM����Ǣl���e���Н;�<�����{�0�d-�/Tg�Q`I$��{��l%�9�*K)�1����~N�L�����l��)����^7�֏��]
�7�Q�8#'Nb�R���YP�d����<g_F��8���lg5p�ww�gl�;��s�CI_-��L(�e�]���v�T�P¡M=]������iB���Qq�q9gU�ȍ���Օ��7��\E
|i/� �_�Nb�MtH���5T�Q�+��5�_���K�F�K�i�:Aٍ粗F F��;��6�II2,�Np�S�S��@��E˩n���l`���bT����'w	++�jqX(�csb��d����[b����I�"��k�&�,5�<��A��"?��d'##}z�Xz�,�)�I�ï@{��8��Z'��$"n��{�|Co�;��yV:����I�:�³��϶�g	P��4;M,�6��!�j��s�Ž ��7�\�!�v�<�|x���	(ZW�l�3z.Ֆk;
������h�S=q����S�ȁP��O ����44LU��S����Nnj�1���L���L2R�����0ߣ߾��-I�,ڤ�P�Ĕ��+�ݎDĞc��:�)�|���p��d !3�j�r[�́�O-k�(�6��染��Qԍ)�Rq�9,�H��é�o�
I�G�S���`��*G�R����p�<�4����ڵh�b���8Q�6j^s�h$DY�,Dn5�&\F#�ͣ��h�Xv(/���db�9�f�&��8 ,{6p1xH��<�#YE���`��BD��-�lH:��U�9>���fh�hfD�1��&w�܆83�@�k5Y���$��XI�S$�<���`���8�7n�6З˙���7u��b�]:���"5���TQw>�m��j:&a�K�G�&�9�g����R�40�*�f̧����FT[��n�<wJ���0�p��W[��s��Ta�]�����1��0A���Jv����Tk���^�N�X{GI:�J�W�/�^�A)RO(�$��S�p��rܝ���Uh�S�iH��,K�u9�-���mq���B�-���6���sqs|E�q^y-s|zBх�A���`�B��bt����+���mI�e�*�Qp��A�C�`�֓�E!�Lc5�n�n��x�H�e�Z�(��O��4Ã�-,���1~Қ���;FP�s�1����s{&�c�$��U��:)(��<�?�w}:��<d~SF��]gL��~� �Og���0Zm��^�f&K��<��;Y��/�K-7��9VUzQ�)|�|�l�ح�D�U��B
�=��c�\%�
���k�>W-]�e�P�0�C��B�5,	3��D|X���!�#����<�!��T��]�����v���a�`u̼o�a��d��p�!�&��6���/���h`�>nr�!�zV��0�b�X͸�l����;|�����fM��oT�7ĖR�њ�7I#��s�- U�/���ꓓ����òD�v^s$����J���h˜�~����of�QR�(�¢��W.����
�@�ky���g2�Q4�[���b�d���#�O?U��V����}���J|A�6�ג��`�l@$�y����"�5��蘇�������l��&4�gWls�z�D9��'�ƭԠ�i�nG0j����gI��ZL�Ϡ�i��mF�7FT�b�Y��H���GM�~�����F3�*���-w�SmB�rx��H�d����B/q�Ÿ�j�74��5X[��G��nճw��&Uw�Fj\&�U�аW�/ڷ�+��R��ќ<i_��K_1[P��@�6�B!�_&a!QG��{T���5"�u4e�0��Hq�ǔ���+�7���W(�+�+������k.��e����RA�P��τ�H���DOLwC~K�����Y��_j&1�톳�p+������4��B_��N��{��٩�#�Қ�H�t���0���)�2��;�b:	�:���zȷ�Pt++�v��7UJ"%��Nc�JK�/>q�gN [ϙ�XͅfZ先IG�R]k�B/���^�M=5���k�́�{�xI���|�䕣��Ry�#�ֈ7%�O�5˞<�2����wo_Q���5J���Ty@�}$�}^ۉ�\5����%��el'y��
*�;�p�I��8�&X+�?!�����(�t
o����g��]��<T��]{���6A=�tA�p�(w�v��>��Hp�C�dt�\��z�%��1��tR�0�_�h�c�f{�mO.p3�l�A/�(��Hz$�5w�ᷝ*�Gگ�X�H���s|��d���ɍ�,����!�'��i���_+�F�>�H��׆oȨ
?�싓M}]�<_ƴ�9X�G?0+!��rTr��1�CI��nk�}td݃Z�m�@��7z|��+ѳx�S{�M =v�#�����e꫉�\ey��#jXC��f��0u߽�5�ӳo'�L'�}�0����dj�i�����Q͵p���/���� �S����9	5��!''?�x޳3�r{"��uUx"$�`܋�y{�|"/T��@�LKE��[k���3�A~`@���h aC-�j���l\j�g��%��fq� [n�,���sOX| ɢ��7�X�5�`���m����w-d�D�љ�/�G�J{����|?~�n(���+�tU�P}0;�&'*1�4<���5,ѱɶ��O�l��Ҋ��$����K�.���Af[��:����i�#�TbsK��M~�L����b3b���i���g��Q82(���l&��V&�-|>�O�(p )?;C����٘oe�A�A�3��lr^y���KcK��:�R���$�ڣ5�m5�YzgޘHV>��c�˜��8��@~��3Cz��ްľ���c�����2��YoX�I�ٓ�ל~�Đ2��l(�w�r�q�:��)�'a]�e�����f�� %@�1 �q��5��ٮ�9p�i�.���-��m�0wU� �\P�!Q�Sv��#�����t�ϧ/`��I������G)��~P���,������+]�^<��j���y�f~�a2o�#6�R�W���u&ǻ�l�`��n�7���)4�C)�A��j��b
gx}�oIS��o2�}#�	qIݟ��V���c�>q�|���k>";|���=ߖM�rQڇ��a�4\��4<�Rck��缕Bq���`?ٕ��ǙSfÁI!�C�9 o����&����Sξ���}��4��̀V�{v^W��@�����w6"�j��z�8k��w���<�V�Y��5o�L9l�5{9*ջ�V��F�D�F��R��(g���^6�9�0�_p8Ϊ0�
*@���!��Γ��7��\a�s�X�(���n��m�x�Y�N�֥�@P����_,�*�S����ҐRT.W#��̉�C�-R��CXN9t��8F�ņw�E�sxȉ"����/2��^�fL����N\Hh��LƜ��5j*GB�$؇t�Tec�i������2��]��L~��o��y�
T�S�G=��<1UG�\s�����.0|��P,K:
N#���\qy-
a[R,lg1߃���/��-{�U4�U�뉊ޜq[U�8���q�ml�hI>��[45�R�aj��2k��I�Jz%�����+R����Ϟ��/ʺQp_�O �%+/�Η@��M:m�Q�da�қ�W�i�9#.{v������eG��_����*�\<��T8�J&3�a{J�~a��?D�0<�%>7s�F�R�+�*���r@F��3�����.W�&�+�o�#�PY}���E)!�-�N�p8���×��[�^u��j��A�a^|n�||���%�Lˌb��:MNK�&��};�ew�t�~�B,=�-�SG����vq4�H!|E�x��qHa�O�ލ��uMB�B���K�Tٵ�@���3�"�P�ͽ`CWߦ�InS�I�ycߧ����O8�AGlz��Z�v[���~�a��,��������������9�7l��s��q�+��������ƻb�
�����-����z���c�/L��P埚��Y�$s�1�>$�d��p�hñ7����KA����?��Gq�� <�_�<�(��R����8rJA�\�Yc| `�ާG���G��dw벶�9uh鬎\��"vqNp|��-�s�!�9PR�#�b<���K�6��VPk�w���)X"��v��$W�g�"�R`N�E��E����ww�΀��ˣ��:�߽�4Tuf?����t�D�ˀ�&��_�i�cp���5)��
x�����Z ���\��zEBp�X�37y _���ޕK$'D[�T��Y�(0;����þ�r(gx�"��a����C;�/DF%��*���@�RP�?_�bvD��&�a bL7*�]�-�`�So?D�yǒ�s}r���~IF�x)ϨJ/����P������E�B�sl�b�5q�4G�����'�S�rs��k]M$M���6��vADu@f�&i��If�'��C�2�V&��U��X��[f��K�p<�p��@�=�"�[0�,����s��ge"�����y#��ĉ�ۯ3[���S,8=ji�rǌ~����~�c�I���fU%,�Ɏ/Ez��k��υ� ��^�y�m���'G���vG!���O�݆�!-³ѵ#����à�1�+�03��s�ÿ�x���n��,����Ȳ >�>���}����\a����e&�;�gi��+�-��o�}A6MD-lӳ��M�A3�C%��=��\���Q���\?��a���Y���\���Z���їF�i��Y+H�˥��P��1�,@���qTU2��'ז��⫃��/�c�o���J#��
�@�㡨Č�a"gR)�1B*�	7*��\�6���&τ�Oef� h��D�HB>�t�cI��O�� ��
ф��>x�s+I��������ͣ=�Nx
���!��i�����%.���	�_��r;~=����BQ x�DA��rw,�5��Pt?�ʹ<D��aU��{}�`��\Q�7�_�རg�ޗ�q���eH��(����:͙%s��y��܀�߰vR�Wk��ʇ����yX�V���(�*�y�
�_�;�%��7��#e��Hn�����U�����5;{8"-ꆚ��3PȒ��Re�s�K�yxb�a��P �a|�.g#�i�S�/�	��2�Ï$.�y�B�l�l�-��O+=s��*`F�jHO�J��z�\��rI>�����&���J�4^�S��;p�����'����{EW��~�����>	�r��7�d�'����/I�����o"`٭R�du�ƟS%}j������������1��#�� +б���k���'XA�B�� ��|����\���c򰞹7څ��q^��+�O�:���A�Io�,C� ��)
���+3IS3ׂ`M����
l��4G��f�4����˾��HDc4��Ұ>w9���z��{�[Y������qRz�_�-^7��/o'[��^�T��t^��j�UIpWh���gc2<�dl��]ŋWfa����	���6|z�v-�r�ތ�Z,/{[8S��%��:����@z���M�Y���C=�-zF��@�|�@�]�c�W�M�@��Z����]z�}r-K��m7�R�Z�G�D���܈��L8m��i�����8���5����Px��T#��$n&d���DۖIܡ�S@��<����U�"z��p
juPP
����s��{�\Ԫ�dqjMP�j��!tf �����+�C��,b�Cn2��ř��CR����0��W���-k���Zʂ!�w6�˭n�"(�@U���`���~v[�h�R���=\mZ�s��e����[��ӑ�,�����X~XT�l�ci�G	"��F-˧�n>muTb�E��Z�;�|vm��6N�@�U�f��sf,"���c��E�@��뤬d1]��N��ff���o��ט]��� >��E�GO����9U8�0�0���"�rk\@�(3!�v��Y�qĺU��O5;�������[�Oƺ)�W��>������W�>;X�C]�jW����s!�c`����}b�����@~�ɑ���VGi$��)�#� ����/n�m��	7�!�lb_�u���;@M��s�R�؏��{�%�3q,[����p�\BX��U����I�(����!�ի�Ă|��;?��s^��c�B����C��x-�a���̞��eGs��\'V��+�r�G��dc|�{�Dg��{s��e@���vt���+���)�(+���֗��r"�D~�:�vA�^�-�ͮ��u�8�)�bT�VL�G���jS:�j�$;j���$ާjÊ>��Mb������]�d�t��?��C˰��5<�t�
pB���j��o���s���IB�OD�ԩu�X/-*�<!2\��H�����D�Z&S�8Ei���d�tu��:Ě��Nݏ��=o��2"��έ%�$�V'�v�`n�����!��9�����e�~�R�0��ujD��l�8���������yέ��mr��% 0��I��|��8�`�:�PL~�<�v���X;4�:p��T6KU.���ᄎ��vmh�϶A��W�\���(��ڨ�q�^M����I�ۮ$�����ʻD��2L����I���"�a�Ť��#aJ�
�����V*�5vjm����B<�<�ڒ c�q�-�\���!$�=1"I	��}�R:r� |4'�GC�߃P����)8�R�'���4�:�
�j�������&�gԓ|�0/�"�*���U��Tt}1"|<&,����h�=�9��^��B��^����������Kߛ]����JħqCND����o����Q^i8&�����@!i�hR�U���֍_z���N3f��I���k�"���~_!���Avś8^y�`*6T���&jp��s����ʐ�jm��
fm�&/MM��3a�~1p��
m�m���E4)l�v5u��������Ԉ��j��e_�7aiլ��;��XQ�֊G�X\vo7�K��,�SP��~1|6 ��br��fR�&9}���U\X�%bM˔V��FÓu�X�.� ��V�c���������H#~ɞylb�v�^-�Ǥ��N�-W�Z^ ��P:i�/�O���X G~H��6���zꢈ��/�J�W����<	�(���c�ކ�	$L"(��D�+���˿`\��O��,��&�G�ā=�#I'��Z����>��U@�{�X�I�:-���#z��lw���q�s"��)�cČY����i�4�9���i��<U�=tw<:��W��O�{�;i@_� q'ČPg��o[ 
�D��E-���i_�#��'EgI.7���=&�M�������oNb����4 
�6�L�3�V>nY�\lI�b՛��l�0ׄ��oj��a�_�2��V �T�/���1���ú-�S"�U� �Ho��w+|]J��tJ�"�����c�< �-B1�K ����+K���\��J��ǏW�Um%A o�"������a�o������,���4��J4I�z\�s�'o`��xA�d2�+>:��!�xX��Z�Bg�c�=��Ǧp}�#���d���U��=j���,!odY��|�9��/��Cq$�ڻ��3+�f<�Hͩ���6����UC��ӅTr:U9W�8&Q�Bɀ��ń��o��C_��\�w�NZ�#B�P�6f\�?���:����B�����$�Cf�����2,0("�(n�(�!��|����Ao5y��(�'�*u�t����~w$��߂mۡ2C�c	1�,��e����_O��;�9������iJ�П�}I������
�+c�Io�hs%�!r��� 3���#�h��Oҋ\�֦7�=��?~�r�H/��	P���h�1��'�_��晚�-��Pl��5:�%J�׹~�f�
����n��˘*w��<��-����$ک`����Z3�È��������8(��{U�����@����/A%���铮D�����!r|���00`�r2�[Ν�+�*<\��%�4��H4�<$4�G�#�'`�l^ű\198��ހ�?3��h)����vδ�dE��O�@$���V�|!�_�+���e�w�EJ�I}��$�Ht���^��$t�@E>��+x��L��;ޡ�0L��#��(BF�vXߔ�,)�V��7��L0�TZ^/+��y���j!fa��1�F�b��f�����Z���V�1�,>��Mw {P���5�����tW�Q2�[�'���+���Hm�,?R�Y� `��yT{�s�����S=���V��!�t3��1Uh{��)L��ȃ��6�
4�N�z����^m&��n���C�)@�V�k"X@���tS�ཪ������������<�ϣ�q!-��oCx�r�?ars��?��;I�3��@/b?���!v� ����|ůǭ��5��a"5��UsX�nG���M����|���a�."/����6Ĩ�L�(�(��_���m�Rr���O6�����B.Q�V�/��Zi��?�-���đ�rB��w�|x�G�`�_��'�i�L��zz�a`�/F,

��C��V�����LA�	���A�F��=���ׇ�mg|^/A�`؝�(�^��>�#�Y�j�O���2F�^��C�6r�U(�db�ϳ�.�Zf��p¡S*ܵ �ކ"�+*���k>v�Y4IƘ��4/\�$���=�c��2Y���hFv,=��������Ml�h��?���*��2\���~SL�j��ݶs°Z�z��tV�Uu���s�C��D�5�Ö�O�n8g �
��ǈ�(�&:Jt��o��B���.3K��r�}����������@d[��mצ8]p �}{i��	Bk#��K���OP�8!�[g�zs����{G�5]�w͌1e���T�(I��s�7W�̌�=�P�&dDAe)��H�7�e�V�מ�܄�0F��<�etH���>����-\��b�J5����?9^˘�<�y�Y(��eЫHBp�La���(PG�ڋ��H������s����8�BF�7�4���V�Ɣr�E��l�ۖ��=�$C�b�)C<�+{e�)H�w�Ï~/h��"��b3|#���'���r٬HPP^����ܗHO�k6��~���1��]:+k�'q93/1N��y�'���x�P�Y@ṯJ�Ћ�c�e�B��+>"�U��,�v�u�vjB/|\ZN��l��<��d	�;A'��������r������L2�G�\��3w���x�w�E2)�t�#Rt����L�t����+�΋�����l뎦�������S[����C�Z_�v!9$��aX�ƫ��M��AOaIͥIUM����d��IQ���x���낝��#Ց��I���'I��S�Y�İ��l2ކ؆3s�#���(o�)с$|}�l ���K&��#�e,s�\�Q}�Ү�!q˾X�K�H^����&7��O����g ���x��`�@X��;aV��sn�/�ٵۣ�i���m.&~��mc_X�r���V�X[*��'t@TAf� �둞��%����R|x�8�0̖^BIgۖI>�7�͖�;��h�ws��(��>�!�hp;n�&˰�>��ڲ�̺G�NE�{�����g��%�yI����o:;���t ��Z�X��C�8[����T]t�x�>�
>�Q����@�����7�L\�,��(��}u��1�y�l�$�^��=Q�!pnuI7{A8�L~6�OR��1��Q��}�:#�����)G)��i��XI_��G��3Q+α�%Q`|��k�P�����T�:�U����#ɫY� ��v�ts���l! �>�R�~�E�"z��fٶ4��ۋ���Gg���!D��3'al��TNxSUrr�C���?���i�W����6���i�۽��.�[*`t(��`�?�d�F�<��~"�әS�42�+���Z]V�J����.H`��O�����8M-�uJo5?j���O��0�JS�eMy��
�����C��z7X�Oq���,˾�@O��:��Y�B��(ɧ.q���[�xrn���.��cp>�
TO4'n{v���������
�<U)$�F���?���'�|#-\*�#m����96�f�B�_t�魚n�U�JJ9A�Q_�s;P骐B����2}���?+�	
�y�rkг��8AN��G�>n�u�t�".�
������G�?]�PB���7F�]�,�K�mr�$�z�h�RT���^����n~���i�z'�́�F�o�? �렂�B�Y�J�K �JSH�rW��cT� ?:���5So�!
�t �������0͡��.S�Zi��`�퉏qTp�#�z�Y1Xq�k�/���Z���1[Pm7�իC����&"��J�s7w��9^���uM��s�/�4{Mg꿟<�oÑ䞊0�b��z�~�dN�[�zĳ��1��:#h@ց>��N-X�%{ڲ�;Ok�RO�A���<�5>_1#�F�BF�~]0gN̳'�L`���eX#�,��<j���8fe;�?.@��P��p����Ă��8,!/�WLS�f@���4CM����,L���fu��r���>ӽ�x�h�YM�S�0�E���;|;;CV�>|�Og]�-�{m�u^�vp�k�0�8��D�/�t'��VenG��ڈp��l�@�������(���7v��f-���奛,�5(GQ��1���
'$����|��l���z�I��4�;Q����-9�1�S���}>hS(����-�e����Y?u�9���m��ےȒ�� ���um��~��eae��>���t{W~�%%�0��ѲI��|?���r�2-��77�q`0x1�9� �'�sY��yxO�.i������ʹp S���2&5RU"v�`���������?L5I�8��怭���	GۯN���8���h���Liq YP��D��8���xqXL���s�A�v<RqK�7ǦˢC'�S@qPo�8L���3��2�E�a��֭�Z�w��Gk��-�c��;ȥy GE,+^ORŵ���s���&�Cqss� ��wվ�&�*ôN�����o~-�zF���2q������K�<��i�f�;w����`bW-��+�΄?�y�Ԙ&Q�F��a�������lB�ٽd-�iiL��þ���r���E�s]�6����)�a��&�f���P��y%����d��x��=�s{%�h8��~�JDoи��4��NV*[�@Q�g:%�}sHEI�wh��=�j��7 �o	�P���"��@K����qjτ�ϛOη�k����i1	B1u~��=���-�ӻ5�J�D�hy"*D)�����I���"��6i~"Q2T��
]�^H%�2^��Q'�*���{ɸ���>˱��
��BI��M�[b���?��UL/ְ�|i�xg~���w�o�s��jh�K.�C�
�=�����b(/
�P��U_�xh��K��Mi
�1�9@�S\e�2+�$����唃M��Z�]_~��J�[�e�C�����9�s�5��� װ?�y�ౕ(^�����%w�(����!�.��V��}J5���U[�;?���e�nu��<h9x��� $������-�XUp�Xht����xf	��%@]����n�n増�d�� ��j�\z)Y��8�QB�	�A(��3I?�\y%%�Œ�2~�C����^�� թ�"�S��L�~b� �9��2�1��\}����h�M]�i��jiԛUFk3s`g�8[��l��ּ�\r8�-S����巧L��hF��]�+ҕ�~�r�!5q:�O�r��.��I��:�!��'�*�O|n�������I��
��`�=�[�
Ig+*�H��r�{R�������E;�چ���y,?���$E"�]V��bl�NZ�O��"�,�Y�%gy��9G@p����\� ��l8�:�x����-;�b�\�D�-I|s��Ѥ_�|����N^��m�������T{�0=��B5tZ�i���!-ՕȔ��qx��S����A�Y�qj��Qsxʼ| skNP_��㓃d��iR��·�n��*x�պ��|��I%�V�M����aV�D;���z50޽]c�%��!����L.�����'��`v�I���Q��߶Ӡ���;22!<72{x��r���-��$pm�ԙN0s
�����e�k��UT�����B�I%xm�h
��*'��DƝ.�P�� s#TF1{�|��f��u��m�u�%�aG��1t��s����]��WlDk��.&A���2�����祓���F�57��^7l��ɍ�G�p��ֆ9�l�B��I]�*=K9��_
��''g�=��/K{���N��������!L�E�����	���RI�ok�Y�څ�^�q��[�H��7nFy�9����o�װs���i�`+��dՎ�y�����P	0gs�.ƾ5��ѐ���]��7v"̱e${��O�u�ʃ�p�����r{5� 8� ��'��'��mj��[�3m_|���1�w;a�H��C䌑\b"6#�,6����r�{M@F^b�;mFS�9/�&�M)V@4ތ�W)�ܽK��t��_ca�q�q��>3Ov8%�F�5���zkX\�x6��c��!��c�����M��+��X�.&6�;Q"h�O^qǿgܹ�g�@�I�\*z�^wiS�Q� p�I�;�X�.��h����ʨW�
�������g:`�VaD옶LO��M9�O�U�J����]�I�&Ji�9`�){kL:��J��el%ŉ�%[D�yi�O����IE_��1�u�[ą�'���/P����Ih�	<*�3?t ��{�4	�:Rv�j��3G�Qm�}��~�z⁑�S^���/�	���l<�@@�G�>�"��b��w@Λ3�8t��4��K�y��TwF�T�:Y�ϦE�o ����}�#�A�7�ũ
�&�Y\d�3���me��`;�.��CVd�����_����ӏ�4��Cwf�v�sH(���ݺ�1�-��U� &��
y3�z�;C*šG��K�3����"8	�Sj ��Haݏ�h���}�J��蝏&O�;Sw{gQ���N��,����k�I��:�ՆX@;a�,�'?���z�m�� ��+YO�s��j�$5�	���	n3`'�d�� L���;��6ĉB�Th/�R%�."��1�v�`�l��>�,5J��Fm�0�ⳛ���P�������e���܆v��w!��a���q�w�Y>��
L��?7�V��f	�dS�A��,��~	.N���Ҏxn ����%+��$wv7d�󟛹\[�u�k���h�A�Q7(s��T���2�׃�� ��{�Ր�ȟ�%214���Þ�1��u#��7�K�rɰ����Ȅ�*��"�������T�K�kT�\ ��v�K��0Ԙ����M�I��ׇ��7����Y�r5��d��5��?�%�K�u޼-l+����\���_LòÛjmۂD+<Og�, �J/k��"��ͅ��?��(ȋ�8�k�u��Ұ^L��2ϙ�� ٩�[X��.�g��l��'��D:*R~ͭ��I˚�d���-�3�w�[r�N���1��<�*��}]]P<~��\�[O�M�J�
�����7q�~eD��8��Ѕ�-v�W�̏\|hכԲ^�p"������P;���;��V���8ΐ��	U��7Ja��n"9�Z�sߵ�؊b�0��h\E�j��5M�t�����]��"2Q�e��Y�Sĩ�+�s$%A{�^�\w�B��:\�N�Vڇl]`�C��Ǥ'���L��ݻ�|��(�6���s�$:+T�\'��~[��J���B_���w�Q�0{����Ρ�Xӱp��{��M�M�
�E������uy�1�f#��H#3ȩ��*����Jz2��8$�D�W��ɮ����3��Z� h��hG
�s.P�ጋ�?�ֆig�C�)}6ƾm�6T�ve��2�G��@��ʆCӴڛ��a@�H�ܞ@�޷ƴ�[����a�i�L��9�r����*f!^g�~��΢�N�*Z,�Q�B����S��תO L�mR?p�O*l0�	��]�sw���p�k�I�a��ogY�a�wɅȕ�#�Ѱ&X8��F<��h�U��25;ؒ,C������"���O�o,�Q��>6c��Od���o&�����oєU�����yE�1ar������w֘�A%&_^��;�Cs�b͹�����H̀�"��`�Ks��B��d�V���.�nQ��#BU ���~�з����lJg�H�:��U��+W���՛��s([�x��'5��R�	l/4��ż��rD��f�jH���:�:�\�z�P��d�2@G�RA�ä���������~y+G�'U��T]`�#r��Sn߁S�,��2^�r]�.�S�|���'��У�>� l�j�#)��6x�ZM,6ӑl�s}α�Ōz{����&�J�Հ��Mz^_*^�*y���`��)�����?ua`�"�c�Z~�����r��49#��h5�e��o����~A
o��9J��]r+w�wt��6�����bD��K��)��L~���.ƃ��@OY�j	#�J�Cb|_�{��ۼ8�� �9�� 7�L_�5,ì�&b ]Y� �JKנ�Z�_-`y]N*z�b4&�w�z/�m>F�*���u$�bq$�A������%�R"V7� Ǽ)��B>@�<�	�M
~A��E �x@�)��g��6�ݐ�i�r�ݔ2��	d�O�b�N�9�f�p������|�*��cb�B	������}j�+�I�^�U�ށA��9J$[N	!{U�S�P��D?�h��A��-����+5��W���.����#)�r�04U���Bs����j\Zi��M�!Y����C��y�>|n�I�_F�u	ۛq�O;� !7dHdR����%�(_�9�p�J�{Z�P7ӣ�j�ʋ���:,ױ���bS_d��A�X���'���F��
��7H���m�!��^W{��	���=�T��V��S��ܟ�8L�B-��9�0K%��N=���v$�QV���LD=�\$M| ' ���A�&fF�w���>�uQ��8�{d��B+���}`f�YIeG����4v�2M�ؙn���~ �*�`�dz��x��g���di- ̏0�`�q�-�����UK�+��PS'G�0H]��5�p�dz@<[�&�
[N[�8���j�&iߘ��XE/,�z�Sr��a���B���VG��0��b�&T��	�A^F��Y#Y�V�}P����W�¦	����<�6�	Q��ˤ�Sm��Qu�WK��4�8�Ɲ��r��Ƃ���DX�J���c�J�֥h���d��,-��|�ը'6�]����O�uhS}�7��,{�?I1��
e?R�zz�����d2zd��5HE���vP�q3�{�U�LQ=���#���C"�X$YNőwq�Y���K��0v��]Q���圙�O\����R����	�*���|C9��+b�=�R�R�S4�w��0��%�d�t	�B�4@���Q�+��Of�qXv,L&��"�n;�}b��$�+OG~�`��~)���pVg�Y��0>�P�Kv�$�=aOs�Z0�~8c�/z�"�O���l+���p��6��~۹f^Fl3�[�ݍ������'�jc�����Y�R�4l��!�����G�
EOV8�Ϋ1db�<s��+Xۊ�����у]t���Yz��W�l�Y��7��:�H��E9W�ZZ�9(} wdm��t]{(Xa��ҿ:�2!VYz`e_ATr�XkDTr�� �8;\J�h �lh�(�R�e��f����q��S�x���/���m��Eͧ+�6��*��H[{t�`�=�"QUQ��-_1}8�k���O�4�*I���B��2T���ĔJ��� ��y��'4y����gh�񀏐q�(��^S��e�{s�2~|k���w�;�Qy@�bl�Y��cm����x��"��ѐ%�(�[;�������j�T� ��_I���1��eI����i���yj�hd���}%B���jU"-���#��\rP�ؓ��Et�J���-�8��6��'2�9��~�O��� Y�,���:����K �<h���eU>m��j!��`���%.���Ω��a CV��Mk
�{�@.O�0��4�ogH0�6]���S"pL�bTE��2?+lX������8�6�BP�_ �8�3��]X�Y��֕��ݑ�>H�杪��fV�����:�A���l�Q� �����;��)a��*J/3���@��;���hn��2��+y��]}z#0ɩ��A0��ǀ�3�~�6��7\�����]P�t�ՠ���b��B�=��n�t�D ���$���,y����[83'�$���kc������Û�V*�E�z�D6�[D�el�]IJ��Jn������wX�8%�D$3��B�����7*���З��A*��V�rȬ�{/n��:��ÂMBr�
k�7���S`�7'	x�=�M,�@�SK��	�nk��}B
��}���ܟ��1�i�:D�]o?n�7N>�IB��_A:���˘u�#�gEC݁a��1IYg�!�ȭ��ofg�]r^N^�= �u}��>]���^)Z�v@��)"}�i���$��A�n|C���#�~F=}x�iԘqt�t�Rj�Jw=bp�ŰA�M��R#�[�7��>�]��b �c��[����ѐ�`߂&#�h.���J�O�dX�#�j4
�ѯ
�כ/�Y;�f���a�5AcV(�B9��T���!���̨�1��f���S�]�G�1+��'-�\��&��V��h,��L�lCf&[�n�Y�|�C����e 0�	R�OS������~����/bTޏ��wVׅ��p��pٲ����>M���Sm`��0�&���M��Oχ'Y���f�īA�5�`~�H5,E�[/�߶U�V��%�V'�4��ד�*�Q�"�F�6sC����n����t괯y��7UC�" fV ��h���Zۍ��$GG)�u�m��)Q�����O�����_ͱ�4]{p�����X�V�m��]J?rm�o�
�P����`�I�EG�c8�'rZUA�Iqc8��l.%��,�3���vL�O�m3!t��Z���
�&��5V�U�!�8�젓E��D�{��u��Q�x L�I,�V��C별qCϨ�����zN��qZ�7��ύt�!�[��Kʓ���fAP9^���n� �=���1��.t�t�HF����ݬ�hڟ<�bq5ӯ�.Y�����<���2�� �푡���_��8�\v�D�a��A.8�䲂Yx(|�Q��>�G���x��EXE,�tl_�v>��]�	_�9 ���<�`\z�>���)��q��RӼ~�!8�@��X�bi�*Xu��"��R
g)��h���6o�c�gPtv��N(�d�`� �Z5�*N���%U������@u���������{)L�_��T�ۙyF �b�fc�Mw��v�f�U��H ֗��u��  �;=��"y}���ZO��CN.*.���Zh �$��
��Wp�>��l�J<0"�3�s��-cRˑ*6#ˎH�a���U���:u������m�]���6i�+���8_E��s ��N�?��~֣\}q�E��&ģ�)��� ѮF�	8�rV���J���U4^Ж�I��T�� ���A���ti��`�cD��"{�x�}�g(<�G�`�vkm�"!L�ԅ>;C�Z|o���*��)(�����C&�_� ��
����傖eO�`ΰ|�t:�]�`��I�*Ō"Y=�>�������ᦸ~���}$��d��'s�P�S%»(Ԟ��!���t�z���FYeCD$v^�ƅ;�Y�#�Մ��xsnNx�cd"������vDE�0`rs���"�Ey��`�iA��H�����M�W7�FQ��qI����a�񁃃��jF����t���y~H�(��@�e)u��F�'M��)Qi�	�H~Ti�^�xY���gca�׮ld��n�{-�%�����^�S��6���w�;�(�w�A�B� Ti2�a6�Y���o$#�e!����IV��R�}ɹ�ϓ	�ƓX*�.���5 �'��v�0���so��'3(M�be]u���~hy^<�uT�A��}���q���[��X]���H���=��e`ZP��	v�����L<�����R�3��/��\q����gTt�h[��j���3�8 �P�����d�לݨ���#�nx��A����_=���7�Cv��"p�<1.>�ƻ!a �uS��5ǚqv��:x��(@D���K���Z{���DS5i�=@�{ռ�������l�k��4��t��pb��X�!�@����8@�V�3��18��������3c�x�~�8���N]��C��	�t}袖e-Q�䉺՜�Csp����w�y�G��qeYl��R
�\fl�iE]�
�<z2f>�����{����<��?p)��}`%~�V.�?����ۡ��Jo��L�ݜ��P�%��<S�ݍ����ԉ���噳m,�a�b��~��7��5hc����ϸe�
+,u'��K�F>L��2y�����Ԝ-�#����z�P�L@���je�k�����5��i����	W�$.���l[Z�O �-��4�[�/1{A��$�H8����?��w���?#�dE�����������i߈M�.Gy�!!�e��Y
Z��S��c�2�e�k)��\M@�Q��3{�`{I�ӅC��x5�/ݍ�#4{�ڰ\����թ]�ZRu��|�r ӌ�dӽ�`�����6'�������ώ����:��XQ`��?����-���l��䄖�A�%��/݆�3��`��G�C1�����x����dLߋ?�+������*k��.�A�����ڋ�'��!�'�S��� �UH��;.�?����N5>���C\�*�n EM�R�M�܂����s�Q ��'y�}�Ȋ�:����3˽�#i%ǁ�R��&JqA��E1z`F�4'��ܤ'ł���kUT�|��x0b�"�`���t�(W��J�Af1͡�RB�g����ЩuemD�*��n���;%����Ķ=�(v�>�-���uH������s &Z�d.�b`����	|�}w�=����<�齾d�Q�KC�U�[�5'#t,��=Sr�ē����O����F�=�y�WRZ�R%7P(��8q���s�Z�W@����$���܋���p��������2+WǤҦ�:(�ɕ��{0��ޏ$M�3�12l���z�~��!��wf�<+r�;�#��H��q������1hU����J	�9Q��p=��A����GhvL��uw��=n��	�'{P��C��@:�P��}q�YW����?�[e�Z,o�/�ykHO��6��_vN��u@e�T�EєRyV��p	0|�s��B���	sSJ��`�W��Rw�Z|��\�Ŀ?I�m/&=yI��
��o�ԟ���f�I�8׏A�2����x`������"�|WNH�DRU��z��z�YĜfCӒ��e�@RV�ðm����V#]|�.�lL���;�v�v�xq���ė
��<�?+��l�U�ؐ{�����TH$z_��&,�� �/e�9�&i1��#�y�F)��+��B����rn|��1[���r��+-�c��_� 7��ecيP���?�Y1�- ����D�<]�>���G��J�8�����RW>S̉@�*aM���4Ӑ�u�A�_.%c�gW������z� ���92��l�	��y0���!���:Y�,6!Xד�V�(��=�{���#U<�&%���뿰���|���)�3�7a����ɰ���t|��^��̲���K*h]w�ĨbU�6�,�fg���<���� �2���eyާqJ�Ş�.!���A���:q��>�q�Wϩ���D�\pf���{-�ɜ�"Z��3�Fh� p��OZg�,O��:~�p�Yd��6���h�)�w|w����-���̸�|��֟2�5r�X�̓Kdh�{͹�5����[j��b�����<(�>y:|�wWLD�|^A6��n���=օ�7r5#<��/�+���ŢI���&.&��u0�< ��6+�E��*1�\V�{>|ĩG�G�J�g�c��W2÷��pC�f�586��QA3���f�)�7��� �X�z�`[(��E�`v���c��	th�.5$�:&�pi}J��UYz��0
-�Щ8�$�`"����j"��L/͂��n���yn��%֠E�|�Wl)JtȂ�.-��;z��x���X��Xt��Qî��l٬U���n)nL��)Θ�e��!�X�(z�CR���B)6#2�	���E�JLAW��|��H�2��ý�v��� �1t!`j�R��î��h�G\�6�l�أ�s椮����y�˺����|Mp_"̺;�Z�z&iY�1�5/6�f�5�2��3	@�r���5U�1�L|�Gm�FzZ�˲��>����W�4�I���7�$��*T3ǧa��"�s�b@ɧa�C.Ւ�|"�~�Fe�cZ�Y�?�m���pO �n��0lmK�>���3���S��+,-S�����v�\Ct�6^��Jidep�*��i�;Z߻�-�/Ƈ���Sj��o�]d�^`�ƴ��c���xT�P�����Oח��'�
�(B����+~��b�̨y�ٸ�6|3��v12��"�\�高 �]����=�S@b�/o� ��xXǞ7<��X-�̰�9��t�r�g���z.��Zg�����L6 ���1���ʝ���0���>z�<	�A�T��V�����[�1���F���*K�C����:�:��A��Ů��ڍ�ƻ֣r�rM���moW�N���q�Dp���,���S��6�^��c:Mu�u����ٳ�)����&����g[� ��:w����<j߀��E���6Yw��w�_�:�m*�aMcZ�x�я����$��T����EL{���}�ǖN躰�~��|NZ�pZᐔ��27c��݁��f��J[�Ac�Dϵ�"v����SS����h�C�釈z�ڗ4������K�S��o��!��In�u9���RT3\L���/�n|���>ڛ�����h�Q��I���Y!Q/O&k~��2�)�Qp�ښ��^(��\�� 6\��+O��Ia�B�� m��e+�|m_޿j�d�W��
�/���2�kg��JP���j��ъ�_�_�
k�@7׎'�要H��o�O�-��PM&�[W<�`���O�^�����̙�t�Q[�l,I��8��Z�)/�:�/kc'�%)����D�a Q1���%�렴�2�r�Y��o��
%�o�M�k-�I�P\���0GQ���|�jf_�X �Ԥ�P�&��g���[�W�[kS|v|(�Nw�C�\b{k���Y�c�{w��m����#k9���
�7�*vs����0QR�䏰�D|3�@�Y�ί����̩5/ۗˁ�
�¿;{�����S�ݤf;SQ?�#!��ƈ'�t��;�SM������+��DK
������8�����C�4Ϋ���D׎1��u}j��(�#S�a��x �<��2KV���y+;$����������`����=B��4���r&>�tf�+����p�H��ji������oϊ��'�Ã���8|���ϩFL�z/x'ff+s�YR4mF�-@���S	;��e�z���0/C�o�N��_2��bT�J<�5��">nJs�
�`�g�0UW�It��E%�g�23Q��EQw6e�VKM+������Բg_xD��b��.�8:C�Y�*���=���aȜH�;���˒A��W��C8}��m��$��n��m��Sd��+n쉹���(��0�dO��T�;�J�[��ws�-,��3Ԟ/$�;���U"b@�=&��E0�K!I�~a8��Ǆ�����S1���f���>׈[ù��}�(�j74���-XA�OL�L=8������10�O�`I+N�ʷ�.p����:�a�F��1�)qE=�� ���w����bs��;�k_F�2��
FFr�2�<��'q����]�����udd�VY�����\��$��G��cht�o��'#�}�GG%��.�xXc�x'2��/M
��m35mr��H���P蠯�����d����?
�˳�ЫGx(ǅ|#��d�5��@�.Йc�#:���0=��o�+b�,]_��_���7�K�Vm���_ ������I��7N"!20ώc��Z#�ғ�u?�Y7�7A�T�<P�Zw0���iV	���:V=FUwgֺqn��[Ў��k�{ʅ/z���E�hp�E@�Ut�{�Q�%�"
7:�z��Q�9 `l��Ɂ�[�;[o��48�;��������O!n�$2C_���
��O`b{��'r<�w.�Jx�U�I�QY���^[0�Ǹ������HVpA��7��mdt���Z[��o�ZU�2>J�h�ýB#�6�~î�u�=��~{<b�����;�, �M��ʽ3r=o�����]�,cf�q(��V��a9�bÖHo�/*oG-�3v���ރo�Q�����zxVv���+����O���ڊ��>���Tm�\e�x73c�5a�~W�*�؎*�7 �;��jU3	`Bs��K�G�64�t����"u\i6�'�A[��p����4�4>�@(�Ӝ��^�J��f0��2yA:8d`*v���?/���t"U�Yo�����F^S�*0��,���!�4�r?�[>��U�֬9C�B%�A�d���֠S�F�	τ0�Y&�oZ-�p �.����1W��b�N\P7w:�7u����r3)����6�a��z]�8ҹ�8����u,m�����`�����ܭ��tk�C�"���5�i*� �Xt&�^�,�׊Ͳ�g�f�x���쁄N�c�uA�-���Ւ(~�|��I�$���h~��r�z:I]ʰ�V�\�&�&�����a�f���%�32���MJh���K��Imv�,'���)����ײ<�`�@k@�Ogi�icw����~��]� �x��TR�����'^�	�ͽ�Ut����`w�
��T,x:`L����s �Ʀ+�C��Gw�,�B���5Oͩ
N;���щ4�B���y������V��!q{�(�<��=�͌1<K�B�>3�/���ڔ�	`�)��Ov9�Y��+�m��rcgpC0%'Qp�}�禍B�����!�\��1���w����^����k
��o����#^�$0'Sڇ���i)]*&r�&
��\b&��qr�p6�t�D���1��U�]�i��*��n*�|Lu�rK��¢�Q��վ�D=���5$�7@ͺa��|:�7-O��|�[o�#����>��ݴ�޻m�>�I__5�kTD��3AΕ|t��X�,؍\���Lf~c#F����<�*lL���"���`-�ᐨI�q+/�kd�D�$��3�>BaFLؾ���1 G�	-�����gZc�-���7O��f��� ���}����]��!'>b�C,ѝ�']��ɋ7���Jw����ZN@U��(�F	�mѤ��ˆ��>p�hȳ�I�s�3��{c�Z�vt��ط��C�G�݋�8�^X%Ciڀ���kW	F<sl}���UJ�3W�ί/|@��l�&G)F[������9�Q+�}j&_.�#�$�����~D@�Z_M���c�� ��Xs����n�k�A���K��秄��;"���Z{��iK�5.�Xc��7z��L��J�<d��x��^oM��&ERdS�ʙ�AiW��D����,��v��aS��\�u�[��<�=��Z��!g�ǲ�cd���W��>�$r�b�?P�H
Dsu�j���'{�z��/���ŢL��C�c������r?�p����NO�� 
�S 3<2�5�g���Բ+�g��;����k_��V���g��xf���O��jjx6vk
٫�!$6�e� *�����<��[��r�49�Q�@lB߬
M�G��8�@
Q��x銫��q��qΠ�7�AK����J�nN~���L�@�'��	�8�Ƈ$e�;�
y ]�{*Zmf(����Za|��ۅ�'�w�k�|0.y�/������-�@�4� ��R<3ط��V��!�Q�l\�Y���|�@2f�Wé0o�QN3��`2��P]#^:Q/l��$����M+ŷ�N�c?��8�?������uE�	)iP얪�j�����eD�K�m�l�/p�V���dQ�h�i�y�-��~�'pi�w,/�G�[�X4>�X���`��+����瓃�����s=5�k��K)-�	��Qւ�.�>� �Z��ݭ�6g�)k7q�K�#JFsQ��`'��Ȩ�)1����v��13��q�j\2F�{��I��x/��ԙ*�'ə~�����Cq�=}O�//vn)8%9�٠EGM�x� ���S�}#q�ePi��W�R��mPPF��r�bn/�S���#����k�i�O@
�$dE��I�bϘ
E��D~��1v��������_�2}�]�����~I���ϩ�-RY��~�-�sP�hDƨ���ԱL ���K�
�%�� /}#u�N{�nvc�0���4L.9�R�T��tkQ�1�_ZǼ��79�i)��=A�Q,M�|�w]�U�v&���I �g��P�F�HS����cL�����1i��<^�&�r��L1L��	,Շj
�le g�K��1y%�,�,��S����Wv��C�?t��]L�f���!x�rn~���_�=	��%Ѫ�������Q��,F�Mz�X,;Pw���/�.6_��4�5Y;���+%��m;��,�.+��<@l{�im��n}Z�Q��k�#��?M���������-d׀�48�G/� y�0�	�"�U
=M[`	�O�~kE��;g�}&q��k<c��ڮn��Q)1BO\8x�9�&%^r!�v���{����Kt6TJ��2#�5�!��P�<W��-�N�B��C�;��/*{)�ܫ�:};�W��+�zw���}Wgm֧��M&Ti/����ZR��ùMn�n�Ivq-*"��5 ��M��q��l�	5^�����\��	����'7��@,[.�~>$qٝ�@���bX?������/<����YR[h ʷX�|0hN�LFp��?�@|�
���4�MN�}ʷ�4mQM��p4!y���2{�]��fu){�zV�v1d	��ԣ�q�
���IK�D0��z$z��Ag��^n�9n���95A�n ���_�TZfB���3���}���d��ӱ�gk�
!@wi�jp\�W*����2ǲV���/�()A߶�Q�r�0/*�Fw{wQ�L�����n5��Z>Th@Tr��a߃��Vt.�)}��%��f�hm�E�{���,��5��f��1��p��1�l��(���-,,�\���!��g���<�?��3�ğE�~�0*�XL}�a�{쓢{-jG�A�$bM6	ַD�"�N�;j9�TS���U:���Π鏇�{ݺ<����Q��-�D��G���D�l��4�m�vi�����ʈs:�=Kq�h�ǅ�{�P�i���P��,��:�gk=�|a�\N�P�f�Ye��G���4)���ύ6BmK%Z��<^��<�=���C8K�p9�G�{�l�'LZ H7����ψ�l�[�))QfB�è!���0?eAHߣ`v���E�c��w��jP��}�09ځН��
%��Ks��-e�U\v1��8�J���N"z�}
�t-��V�9��T�4g�`���UG-5�N�G[�_3%L�I-��~���Y��t���T�3[��Rv��a���r��O�=�s�����@|�<��<�3�R�$�Xɶݒd5ܐC]��i���צ�`�����>���js͉C��(Ė2V�#[Kb���f�7�.�L�Z5�L��|�k=`D�(Z�A�ё��I�R�S�BW�]AjR���T���@g툊�0>��ZX�~<*G�S҅PF�ɘ���َ��>���q�7��A�QUk3��#Byɘ��H���^WPpFK"���ߝ�+����j?<O���Ơ\h>�qH��Z��&��e���εkx:������jw�
�LB`~~��q���_?�N�nc;�So�FȘ&����DI�8@؋��͸��<o���9�sQ��M�&r���^��~%��Za�Q�|�[D�lf�0�P�1����{B*��yZYe��}�|p�����(��/�g�=��BN�r�������&�1}ܐX���QR��J��&�ot?7C�+�H���]��f�s�Ĕn	 ��wE���9\�_!��9�ˋ��(�n��-n��)�~�X��6R��-S�L��]��:��qM�T��M��dO�R����b'O�:&mt�D�,:��R9�t>�hla��¾ό4���#���	�什 Жr0g��������iF
kƩ���2�µ��SXC#�~0�	Ni���؜�N96o6�V��<��.��e�)���k�-&�U�iA���{�������*����YI
���lA�Cb���h�?ߏ�����qD��lh$洋0�:�/Z��ڎ%��`;��6��ij��i�}��~�K ���6� ���*G=Ƅw�m~���@>���L��$�`� L>zl/v+��\�>�n+{l�-5��Q�*�Lx ?#��}-�t,�n��%Ռ#a����7~�w��QE�)}�1s@t���s�ҡq���3��i����K�Bæ�gb���b��Q�)B���s-��g�Q("a>4�z�Nץ��gG�2�jq5�|�cȄ�K�t�<7K�H^��'�D��w]��>������=1�+���M"�����Җ}���id[q� ��b��Y޿Y�ʆ ?��&�y�?���\w
��$�a��� �$c�1V��=�6ך�/�)�[R8��O_,Qf� �֓��1���d�x�]�w���2��8[�W4b�D�˃,%Dc�����76N�vn/�G��(�Q���uw�,�f�Ȍ���P�{kP�D�8Y)3�@B����unɠ#�Ǫv�n�O�+48��g�*��K��n�_DvS2{��4�MMܘ\%b�$�I�
��|�ǽi;=_��wy\T���G鮭���q$A�'ȢL������� �"�DQb�opD�д�����Wx�u8b8 3�J¹��/%�x�-���s�܀tA6 �R���ū�Wܬ��}I�� kOaƽ�/f`[5�P�B#�ϱ4�O��ii�9�3i�d��甒}K�7�릇��`��_i�B�>�K��T�3I�s=$��(���k�J�l*4���l-�'.���ڍ.�dN�����qzl����!�J���`����Z������qs���~����ھGw��؊�͔�W$�q�@��!�b������@�	y؝</��D�ŉ�{8���`����ql)�q*
�1�nضu����˱p6C�<m�8N�c���Qos3K�*��z�c�sx���+��M�)�fl��L*��fA��'娛����+9��9a��G�����;��.&���S~��fF]�ͦ\�e�%�3�^f��=w�c������V����w����FV���<,�	���1�(�|֦�+Ƽ�=U�S�
]҃���t񎪨+9a*��ͤ����⓯��Օ�a���aL;!Q��r�e��Y���c�ab�^�=�姇 �pxg7a1��a����=�Fy`{7+�K�ps��Ѹj�Z���������b�Z�J{8�ܘ#	o�O�OQk�1��T�x[�л�Kr+z֏�-Eol�U�����0���$��7�
sA(A
~E�Tz^�0��l�_^�4�5V�op"���}X��d����3Ǵ<ؚ�H`0Ě+@��Z��gf�_�G�l���2~��O<���1������Ӗҋ��&��0K�	����}<'0�Q�א,7T�}=�k�R �aZ�n� �[ל"Q�}�1�m��?q�xI$+�`69�z�-���h����A�@����,5���L����W�����N�O�)5�n��TA<@Q������O���`eX�����ǘ������H\����L�� ����F����7��İOxu�0�P>zO&���I�5-u���5)B2=/B�Ŝ��>�ua�i'�DSܔ�����)��FH��l}��sT:�ͼB�dwY�R��
t �7EZ,�6G'w��H�\Kg��4#~	n�ңZ���T��l����ې�;|���Q��H��:���eg@��/�^&��H^al;43V*���wt!_�w�CiR("M���X���ٴ�͔q2��Q*G7�g� "����N�t��u5J�Asܜ�,W1�˵p�v]լcЭ`����RW�/@��X�u�'�8<����-<�^�����0����`;ש��e3�r���K���NNem{�!\p+�%�mE�D&
����'���lC.��d������̠�}y��etW���O�ū�d���{S���S�P�C�ċٳzV��<K�ϙ�/�
�OȓV����h�H��}��+ .6��4dF��T��P��kP��>_����y�=Y@��Ŷ�y٥�hf���oQ8����:���]����ςCA�Z?��h���2����<�\��ʱ��RBo�/sz����v�8�U��-Y�CwÇq�*\��a%LSa���2w�.J9���o���/���z�%�I�� �d�9E7����w{[��[��3�e�$j����@y.�ݏ�:ҳ���	�٬h�~�#x�{a��Bu���	"z�g#W
���d�/�"�� |�*-`���*@�F��]��b�P�����f�?��.���ۑ'�j6�Vu7(�Sm�Kj��X��s�x[4y8[�1��Ŝv����������=z�o0ʟ��?=2�m:��l����կE�t޲9Ψo���V�xTQU������x���L���k��z7�
Cs��.��_��)^ss�p���G�k\m���a��70ᅿ[:ڿ��NT薿q �i��o0{�n�6�y�\�ބn�"4�@wa:���q�*�N�+��\!�-Qr�5;yif�d���c@R2�M���{p3�l�z�S����[+��Ǚ�\eX}�6H~��R�!m�a��*F,V�(���Ucr���D@�%�v"��?]���ڡ"��o�{0���PN�C��$k�`��B�r���b������!\B	�on o�q�������3��IdB�q�& �L�/29�o��~W����GH�A:��]C���ao,�iG�7���
1�q�9
����U�u��8n
�J��ݦt(���k\YC�Y��f��sr�b���C�x$�й�R	��qKM�h�~�x������`��-�
�F�^��w	�T�¼�ai�nX_�>m�M�i��c.R/[�.;O�U���AHd�_M��Nk=�����p�9я�,���>]�5-�(�7D��іr��@a�F��5	���W�棱)�~�s��?S���T�^�%�Q
"�)E.�
j��!b1ʩ���,���8F}\Hi�����
��O���!�������@�Te��m��B�[����A2��*�>+����O�d����+"����������:��W�'���4�E��Oۑ�)芕�_�tĨ������i-�v��Tc:w�.T�+b�3`k��j��s��Nǵȕ��_��%������߄���JQ&�F,/z�ޭ�	-ط��T~�����^OTڇ��}�.�v�))G����qF����.a�_�aEi�#ϩ; �:(�Q��$�5h9�Q�N������Y��W���xr�rw����hJٜ��j��Hul�~,��Å�fo�Sb��A���F���6!���m����G�m��i��a+a�<�N(N�~Q�M�Dr<�Z���l�y'�AA#B��@MGYw �[���0�<��|�c{͠�>^G��)�c��0�b�x3n����_,���Uv�h��̱����B�����b%|O	lE��ݻ� &���P�������H��D��WȺ8��(8`�$�o�8�&�Fl��nx�*m'i�*jش���ɔk��ѱ�6 �';%9��ep꧃���͗A"_��f��֧��h��F��'�}����5��{��v���'���IB��~_�����%�� �����Ncp�v(�{���$�䩊�)1}��S9��W���p2F��W+�M-�/���F�����i��F�^HYÝ� ��J�C"��a�f��E�*�&|�bO�L��J,�߭���%�.p�Z� �@�L�[�*�t]�k���� �ҕ���ٗi����υ0�ɷ�	Rj\��Մ�����΅��?�+�c�Sv�؍��Y��$Xv��_�:G�!�`3D"��d��ڽ/�Sm��[=;5�����X�U-��DQ�=HK<Z�z�1�jRT�[2�Ճ��D�=Xv��b��E��Z8�@�?�r�-Ե����Y�O�3���h�ҿ�2����d�{��� 1����&S�!\i�N�^@y;����껫��JI~�p0GP���o�v�|�c ˗+�X�;��o�V'�B�l9��t4%�%`$E��&4�fcv|�����T�����[�a}��t �����F���̮f5�h5r���d���Uƞ0k���+
m�x�eNt 1>�\G�^0��˄a�<��A��v[�|�P$Z�͹GJ���y^'���'A�}=�1z�&��Zݔ��aS�}=�[*t�����X��>@�88����S�I�c�	Wo��uR�(r��/��u��zj�O2�g�z��<]�<�c4�J��;͊�7��s�0��!\P�O�W�_C>��.�#;X�R�,p$F�a����mC٣f鄙�W���.�n���A��Y7,Г��X��E ���')�$8H>3�T���Syg\����6>��z03��_v��<��_����A������D��B=boq�v��Ƈ7����y�+7|l�	��
���m�T��F���:�����٢8>�|<�vG�+wD��%vkN�3�؊'�)���/�O�܏��I:ę�@�v�@:
!{������3�y:3�X�2zr�#�j:ަ���Jw2��3��S������-yKʹ�;u�K)�����4�,䑯�44m��z?@�?(
�������A���.��m	�Y�NO���ZC����ٵ+鲚1��)�FC-�|eO���M H�G /H��͟�zpgY����_P���U�5a�p�}Αčiİe��a��h�O�'����������bx)�G>Fy��c�uM-��p�b_�a�76��hӫ��M߲���c.Aħ��-Ǒ�80��+��zݞ��3��o�r��B���r�B[-P��厠�v=}Q��R��5"R����VK7�����]��.���RHS��6}����rk����j�o���O��,����(���-�e_61	q��\V�&"�ˏJ�N�Y�!�e𤟛�fzh�6�'َ�Ȉ�����$�,k�W>�U?e�{{���
"�+���h�r����@_����:��'ʃ��<�t%��8�E�v��Mm,���,|#�(g_5��O���!'g\�i�n�	[ړ��H]�]���%��Xvz���̄���,J9T.�/~wU�������okWqN�aM2E=�ֆ��1�����\e3�1CP�V���vgw;�ϖL0�����ݲ�?������&��d�oL�/�v{R�X���"k�;��e����f<�e�zH���G����y��P��t��n���x��6��n�� WX����7�c�����7k�����|��7����.D<��7f�_���	�2c����c�sB�B��:�� �.b�;�e]��T3.�ĉ@��=Mƛr�+ULL �.^�!WGP�@��=���2U���*b\�#TMw�q���~�ua�P��b=�Ǝ��J�Ǫ�}���́ d��TC���DW���Ǳp�)\���Tڕ�݈Y�ц�J���R^ܐQ*Ήp
[���!�?qZG/9t�v#�K?�9p�Y��yC��
���^E9��
4#��W�|}n��M-����˼�S���l��o��	B*�&��{�&�uT�����B�B|3H�h����;g_�� �+��������dI�b����͙�jٽ��z� ��  �t*Ӎ�Ro�!�žn��b����:�r�\D>�@z6�.�X?���a�Z�N��5~.P���"'���~��s�
mx%v2($� 4�S�詂hH���g�Y��w��h�&��upm��y����շҘig:"����JJ�9�v<�� �;	 �}��B�A�)���To�Y�g�/Q�d�����{�ӶyX���:�㹉e)��_��f��)_�A�s�5���Ӡ�ă���QbC�V,�o�5[sL�mH�����X�Q�E` Z�@�L(���;t���C�W��7q� qB�Þ��Q��� Uǝ�4-�ɖGl�d��C���-��l@<�B�QvwS��]��"�:Ѝ�����������3�2uXZV;⼝b`T3{���A�i� '�(�=��]��B�P�[+�V�ܝb�^��	��=��q@��I$Lj�h/b._��J;�QՎ��$aQyI����>s[Tp�D2%��6�b���.�aM8uEa��r�xx�T�f���j�,�Dܣ�FΏ�2U����9��F��$+e
q���G�����=K����N����yM�Ϧ����Ay?�.h��:�Rl��XN*M|���+,�ד�����d,��:9Wa�� ��`V:m+]E��C������j�:q	�Q�1���@U����<��޽i)8w��i����Q����g�D�n�ھ2|��I�;F+rI�,�q�v)��v���'z���lG.��>QǏ}#D [��9�����K�>�YI�����2RE4��7��8�,�>c(d�{^&�(!����7�Sl���T��; q(O�Ͷ�o��i^��c�%Ν\k4�'{O�ޤ0��+�?!���l�AD6=����fne�\���f�s��M�׃�@�|p#�R��y��kF�Ck�H�/�B����}��
tk�y��CUJ��J��ܔ�/ XdI�ug�z+���:��?���i`��%��!�-��0Ȕ&�w��)�8��㍻>����mQ�w��%���i���Z��j�F�aM���hd*�Х�� �@��Ϟ¯�w|E-���r�×��������(!h�@�e'
��^!+��M����T�oU���a�oN�i�l�=�oD��������v6,w]��K�4@�}�A���9�r�j���c�n� c��7�栐CB����Ƭw ����NWc-a�:��N���1����B݂�,����P`����f�s	]��91�^js=52,�l8�A����Y�j��Г��bC�z3���\�+�(�l4��-Cr�dږk�W7&��l*�MA>k|"_��[��Po���!Z�/,�x�*�6���@ s�v�i`��H�"2Z����(�����Y �&l<[%u7X���@��XzL�� �鎄+Y�m�ы�����T���[�D �`*%�ݥ��Q��)��ꇾ�K,m� ��"��q�z4�X��p���0K߈�3
�P>B�/n;��m��k(����;�$/.w�wq�*�oB,�Յ5�Zb!xJ��ۺ�hA/������q�W}A�����Z��`���t��l&�7���;q��݀�?�G���S�����C�������$�Fv�
���pyTh4K[� �6��o Ӳն��z�8�ӝ�'D��:e�|���`0�+^H���7����YB#�8�&�=U�:6���QT׾~xkU�j,g��_�8+����zH��8�YB)�
tQ�m����<O������.0�jD�'E��?��:a(r�#Ђ��3�s4���wv�wMZ�\gy�Y�*EP��y�2m�dj1zR�܏���~5zw!�u���m��K���
4[r��3p���"O�wC�?"^��1� X�͜��h���L/XI�~�@ό�M��d3-������xđ�����fN�.�g���a$P��,���1��ĿB�Dǉ���R��c�J<z.��k;A}DX��F��B�MX��b�kO���˜d�"H��Ys��k��p��m3W�T�b^AX]�I�&l�; ��&�+�F�H��w;y>M�4i�.=�C�ŃO�������o��P����?O���ϻ3�G�u9�R'���Y]��u��pA��r�
�^u��P��
���F|�cq ��n36?�ӭ�,Ѭrm <��^�13*YJP�p\��#= K�����l��@؋���PTY|�[�����:���~����4D�r\q��yo����D����)�z�=1J��ShC�Ej �3-�� Q;�дji%_CS��B��;ؑ��O	1;&89�����{d2�ލ�n������>�D��ռ�^�� ��o
�E�!W���K��L�����.T�n����?��Ь�G3*�6\S�`G�ѽ`�����T0(�˘iI���l�.Xwro�
Rw�p9�Z����7Tvh�Ce���0� H	��D�gZ8E��J0D�ƚ,܍6��׉��U�#4�X0K~n`��Y��?�;6�4�k��@E5ug��B*�f�h@�d���^�P�Z((<f%�+64�����H�Ru_�'S!��>�u�A��Bg����M�9w�T�6���Ɖ�W�{Q��xQ��M o�g��dF�hID��p5j��<)%�X�r�	�����Q�"�/�W����*=��s���Q��q�Gcx).�JcO)��jfo�^��A)�i_X�;"���-s�׊�_�06wM�p�AA�&�KR@�f�j��8*��v�����q��,�/�XP�z���?� �	[����6U��RmGp@�APkf<�ĺ5PzJ���[��ڗ2 "�̀��ch�f䨧��^���qi"��>LgY_�(��n��j����"ұ.[��13�0ԝ-�ZVzz�����oL�2�5�䣵y� F�#����:�}Q���'Y�NWx4��tWt�MK e�^J�f�����J������篂@g���m����%Z�6Sc=2ΖP`�њm59w���gma4�x��y��:Y5�5���`Rk/�`����4����y���@ ��RU�8�'�xՂ	�P���iGm9j_;��D7�\�ܔ�j"� ��DW#���C��Ck��ߵ�H"ﾛ�A&R�B��hd���EW��rc��7���*>�hZO �M������<2#�����2��w���(A�m����L���7UB�aѵ�P�{�Uq�/5�M�����+,H��Q�U�1���΀ƍ����_�޴
ɕ*k�N��r�q��h��\;��'����&��CH)�M6¬�\VVa?f����F�A���l�ٺ�'��y��4�f�/�NH�?���H< �Fh�/|�b��N�ٚ&]�iu�-�l����2��}(m��w�6G�;!�t
,e �A[�a���L����
@hSn�~އ�o�z���8�+�lu��n�ú_<�2���=l9|�T��8K��~`J���M^�u]���@z���a���x#!80���RG�~��������Tֺ�;�$?kɏ�
�_K�l��݉�(�Z��z��8���S�f�����RZ��Ll[vf��yiA���{]BV��
�j�5<�AJy8Ȁ�����`�}�~m�^>��*m2H�|�J/�w�R�MW^C{��d\�a�)�����M��L;�#���+��q�E,䛓��;^J���5��ǈd	־/?��N����Ƨ�^(��$z+��@5��Q��<���w;,L,�����M~^�w���M^F�,~`#�ݞ^��VY�S;���z���O܉gE��a�K5��������P���qE�� 
��*DՅ3(�'�P��xU���a�hrR�`v��&pZ�^d�|��i%�&����w�-������O��������c�����Na���NդXN�v	��ǿ��
`��q���@�UdY��츴��〄��8� �^d����z�Gҵ�f�,��FD�G-�)�wv7�[mj���X_�e�I,�a��<��-����On�m�9�9�Ѵ�=�m�l{cS\F���R�B<2�x�bC��r�/�a�L���ʼ�Lq_r�/ �)o_&�0�:6�]h�K�ҡ�j�hV��f
#?�k�����\sm'��.~�~YG C<���v����x�&�w��E8��������*#��ڷc��h%��G׊M ; ST�Щ+���k�8�ٽ����x���n]�׉��m�ya&R>��&�]M�w�V�B_pߠ��?L��T�E�N�6�Rz�hԃ�rθʃ��H����Z� RH��r�!i3$���S��{�Y��'95˴�Z�P��j|�z[�*Z��2%7��;B�ZX�\�{#ʻg4T��2x��ā�Ɵ�g�Z�oF�l4�)�� ��|Fd���y2{��1��e$W�ƀ�fڀ<����
 4�@�������
Q�Y�U��ёa��N��4	��8qmJ��eej�����'T0t�ߢp��<�7W$݈��L�DW�|�/��w�"PB
�8���ݹ����'ۓ.�7o�7����]��֠�UhxJ4�K��Ĕb�P$�����@Y��}��O*]M�՞��$���p>H�ڔ��]�7|8��t���+{K��w(�z��=�.ʅ��R����$ =���3+�>�х���U�g��<3� =kL����&i �ǭ�x�B����G/^�H2}T�K��X��oq��ٮ�*p11h��|������6�ǊS���j�G�0�;���h d�~�x;u�Eyןq�j�Ni��r��El�%�D*ڞD�#(�]�@�
�\����1
��z�!��b��趔ш���L����ظ)Ӆ=^�w����j�Pst���&B��M�T;�s+M�F�)�oX�o2�OgO>��r�e�G�{�+&K��W�B�ʁ� ���v������pľX����m��Y�c�p[�OΆ��S���Oi��M�o$֋i�d��ѷvp�KT	qHO�;ҷw��0�p4��y�X�{����<M��#�r�O֘ ��UN��{y��8c���u��(��6i����^gV�E8�$��]����Hk�,^���������yϿ�h�7�H���ȑ��R'�� �n�ӡ6iW U��=>s���݉�d���j��; �ic���8n㮼S8\
���c&��	�_���X����ԣ��e4d��6�*w�i �x�y;��!M�Z��)n���/��y� 96A������L,5��+M����+d�B��ٌi��5Wd8�E���{�,��oy�L�@׵fz��jf�Q�������<0'<�|�-�����Ъ� i�P��Z�M�h��۶y_��Ea~Y�t�I,��M��e!ts��*���$A�.8vv��U�10�} �_��L6ET9x<��R�ܑmϪ4�M[4Lz��#>GS~�m�[0M<�!�#2��0�RpǏ��U�[�nk��x����?'��Ʀ��ȑa�Q��e�ko.��I�h��A��0�|�q�F<�W0�E���;�CՀ:�vhޣ�N����ׂs%�̖��=?���iT�ݢ|�pl�z��>��͐���]��=1�����?r*��''AG�����-��|� ����~�m*"�LLrz�!���d���*�0?�1)��n�;������hKS�U�4�j�Y�� �V���I�G��������oю���,uٗ�P�K?lUz�Q)]։�f��D�#�8	tc'ƋNj�݊�� p�~��&�R{)n�����;'���D�;Kgh�JG��uz0Ƅ�7�Q3_;���?)����:]�,��C�L��+�Z�{,ג�]�)��4���^�!�$aȴ�˕�:�D�^!��1JРh�;���R����1�wmh�|0u����9`�����'��O?�ϭ/���Λ"�����-C��r/�c��<�_�<vщ�8�u!Hۀм�\؂X�����|�W\�/��n��ۭ�1��9�g�Z#L��(��I����?��Kf�[ݧ"J|����7{�uh%�[��]��3���&��7H�{�#��x�]� ZӋZS��XM��u�=)�y�I��1k��Rk��'K/�Vñ��8�$D�xO��>�l�Cۖ�)G�t*>X���qF_�I>Ti3FP�+���B����N�uZI0�w�" zC#�9��x�[��,Rt�J����ȔyG����i�w:-t � ]�C)�ңX�	c�W�0n"��m}X_4�W�jcھfh��������]vs��}��˟����X�eq;����Z�Z_� �~Hqy�"�T�H�����9�=�Q�4�^Ny8R�?���or{ ���'��u���Y��ƣ);,��rN�d�(�V\���zsQp��Ɔ^���Z���y��e�=6�,�@ �u_�ğ�$�,J����Go�wo���-��A�t����+δ���-������J٦�L�.�,0f�N�X�fY����P�F�C;��n�B�#�O̓��qLY�BZ�?��L���k�І�ǃ�Ӄ��׋c��Sպ�M�ǡ� ��x�wz�����]bV�ޫ�QbZٰ�}v��@_a9����!��¸�ꦣb���%�S����5�<T��Bߒj8UD�!,�qzf�X�ԥ	3�}��t�c��Xt6Un���[��~�4��ҋ��4t'K�|ͳ81�h�*ɰ)�9��Y;�@1���c!�H���i(�6������nu�ݗ��Be�'3����N�2g�H6VG��ZEp]am쪩@�0]�%.J��q���6k���\@S:�YWi�~.������C�����Ո��t,]^ˈ"Ͽ��0ۑ�w`�[�]�_�/r�����hh`/_q��bc�9E��7�b9y~8�v'���ځl�!(R��mH�M��OU ��9?�'O���0|�u0*f�ǒ������������o4/�?��E�EH����<f�;(��/���B�'(�
�	eY���4:����7���i�Ǟ���j����#�?P����g��i<p�Q]w���uf����0c�n��ěQc��BH�tb��ys��
���6���,�wl�WyoX���m�HP,�q\��/~��㏤�]C:iO�e��c�V�AF�KD��ree��h1��~vGQ*Wй��>�_�-�S��ȶ@�P��)w�QCKǗ!0U�B���]Edk�'�0 ��#2�Ù˿|��䛓�2I�8���BS����J��䛱Q�+��9�(�B_����z<�w8�����D�$x�-���G�P%y�7��z�5��	J�B��8��jtN�r26R>��%o�g!�0p4�+��n1Q/n��bkg(����ԍ{���MO��{�"L���Q�c��b
��;D�)��Ѱ=u�S���=r�xp9��3@0�R�@�ɤJ�7m�p��$�[\ș��ӥ��ۆ""�_��u^Ű���$�T�&�����xx��R`/ټ�}�>�w�x�UV,�%|2�ui�Q�����B=)>��&�X��_�s�S#�d�o�]{�_��Ê?��P��v�C�];ƹ�3έ�VQ�0�s���}��&���Ea���Y<�g�fI� ��⋉V%Î�G��E�ih3�*���͋Wm��/����+ݕ��E"�����ڑ;ٜ^ZɃ�dR�6ʃd��?��qn�c�/�s]V��6�%���6��`	�^�2�D�]F8�h��t"|�ɞ�Oӂ�gh`�r��x�𳌢@f����fuJ�ҋ��2 ���E��c�=y�O��_؝E��+�(x�^�"/����+�O�E̤}�U{����:TNj�v=d7��-V�iY��k_R��[�*N1qvX���p�T[�&�v(��N�2 3в�%KBu w7j)1��*<��\X�%�Q4C:<��b,���y��RN)���|�Y�Ig|���~a�㛊�g;=f����<1�&o�w����%���f�yi!҇�s��E�S���p}F"���GD�3P;w$�˥"|���kɏ(���$2k�Ҽ�����3v�_����]�HOe3M-�2�]�0q��L��g�1\�y?b��b����*)��:^j�N?�LN IރҿI�-��q5Oq6�j�<�m���:�"=����ȭ�b7c��f;Eo���)/�J�|�C�F1E^��A|F>[�Wj����[��?���@�V���̕��
S3�(�pzܩ�wAE'3ׁ�78;�$�V��ҳU6YVu�xKH�;��F���M���˦�u��:=jr�� �u!�Xm��.���$^l��6�JW���bޢ	c�`�����=�ca\��w���m�t`�0]��ޝUK�tp�פ�L ��e���w�Oi�Z�����ю.YXu[O8 y�MُMݍ�es�Y#��b��?���r�l2r��|��bN�^q��G�兀?�n,+�2�qv�8\ZS1��ZfG�)}�������1uhyM0Mxʇu�^�?�b��[����/s�a���ҏ��7	�l!^�~��C����;�(��O�m�hJ�.�QGN�iY3�����[�aq�E	Is.G�h*{�і b���z���$�2d¢r���Y�
����P�g��j
����z� Gp�c����i�?�ςD:'�1��O�^<���mK�K֯й90�����G��Czj� ���1���uH�k��i�dp�׶��(`2���7y��$�er	��geZ�6�:�m��O�%Fy�xT]3l7����'o����13�͡r)tNML�+���PO5tz�x�d���]�{|g����ǲ�U���E�4LK?�JtÑ�Ulٽ�^K�¶�G�� `E�pcwhn��xi3��Hy��Z}!T�th����DB5��jUJ�e�T>� +�!e����y���3����x�`�����g�RW-��bZ�s����[��M���si��W�ek�vZp�Kk&�J��S���{��  ��>�2O�0����	��G(k]U�B��;�Y
<0�L�8��ܒ�q��;�Di��ʙZ}Ʋ�c�:��
����D�p8ȌD�:6Ѹ�k�(	�԰G��T��~��F>%d�+�CX��~�gv���*���;H�1YtY����p��-�Ti9���G��� 9�Y%�h7h�
J�0�.2��E��Ji��k5�v�d��F'K{����ȝ�]uP�i<O^�AC�؅ܠSI)w���.�#@b�AKF�@ʰ�^���w���D)B��D�,pa�G��[����u�F�۫���{��Y�e����&J����7���݇�,��aЃy .��'�)�>o]ٸ��K�{J�(a�웤�Ƀ�,����,һ�u�(��=��D@�0�}QU�N�`���Be'���:�F#�_]3���8ld,�w����K{��;�R�{{��g��e���B=7������=��;,7�ؽWW�K�=�4Z�[����~���QXT�=�������)R��؟�����
�a��f΃��Ė�4�y��1��ʽ5�߶���nn5	�����䣾��~�C��>��>LÂ���M���� 6at9U�^j\�:�Iʒ-Z�K�ܵV���]�U��j��������>�K�6TG���G�^n�/�Se��V��y�)���>NF�&;��PB亚 ����C�b:
�D�Xga`1s��L!����!�����Tq/�7B*O�a`3�'�_#�(��9 �	w�0_�����n��<��

�附$��H��q�9�jn��
���`�.����|{2�HG���n������������"PWX�$8"K��~$)��7:�J.KT��s��nBH��Tj_���a�k�Kz�J�f�Ь�9�g��ɔ;��3��.x>�F��U8f�ް픵�7L`�\j �]��`��d��_���e�1)�H�X	��8��ќ��e���]"es��x�=���}���X��xD������}{���J��D}� �.�,})rA���7M�+���S(�)b#�b��(n/d�����ĵQ!�/1������l�̜�A%SP8���; ��Ɓ��O�r�p��"��o-'��'­��;�Qn>��Bȱ^r�{##����^ j�H=��Y�'縢
�o^+D����u h�٬D��}U)�l����3���1�{*�AԬ����Jk��2m�y�<BP�����ҩf���N뢡��W&TaßJ�(�x�v�S^�f3�đ��$b��T
��r*�&+�Rf�Li�i!��ٱ?Ȇ^����k͎l��.(��1��9��`j�|�Z{8�%�@�nЯ-�
�.R@㉽�ya�=]3�59�Q��,?�`���J�����-�� ���V����߷�K����)�e'��J�m5�T	k'�	�Cz��C<��(p�vLѺ�sBȔ�P=U��5�@)Z�|ʻy"�ɫ~G�[���y\��4Й�y�a}�2��C�Vp
���ѫf����-��	X�&�-���_[Mpq�P
v$���%HاI�g)ǩ%LfY�z�9��G)��6����x\�X�S���ĺ�쀳<�$� c����4��G�DcP�Ի�4�Ӑ���Ǝ叒,5�Vҷi���o��"��r��[�A��j�v������fb�Y�՜�ZB1|$�sP����ny/Ǽ�ǧk��X${� �4�͹8a�ѥ,=.\�������e2��A���W`�y����	�kXPXM��H*S�oR�N��K	��v��A�y�8��Sy��s�gSѕ�%.�y��d"k����#?��H"s��]S�}��E
��L���}>�-��̟ż�M�V��9�a�D�ao\�3qȸwc&UV���7�s�`�����}f��V��R�⁓2\-�f-��(ŝ����kym*r݋�ZX�u��F��?�Ia�t<��y-P �Τ���-'���t�Vo��z�#�p������y����|����}Lp�K"�B�#�c�G����� �~�`֨�2�u��֘�H]��X*ά�����K��s�.r/������wN7��a�' 'P�<P�Pz݋��䇲�WFS�,���0�z�WbBwK`����^A��ňd�5�V���1���O8gA�
d�<Q�j/7�;��/�[.����HU��s�"�Ԩ�ԒĹ@g��<3����8I��f�:��R�k2����rJ�}0�b�VnY�0�k<g�c��gF���P�	��p6�W�洓�>|-��4��ơ�e����e��8YE��K6��X[8G�l�`	�����j�S���,$4W,�W�ĉ0=H�j$���m�*�(w�Z��kA7:�qF!1�ܝ�:�����t�Mhn������䑬I���$���Q��1�ɚ=Z��v��θ�Tyb"���k��cqh�Y+���7�z���I�;�N|+��K��U��w����ym�1���L8��i������80ڑ�'@����eRM��`�9�ua>��bAmk���E����<^E�m�P����������XZc�]Ώ(6+W̎��;����x�7N}��W-T;�6X��Ȅ�g�3r�4����S�w���r��F���`˓�o7r�]�8��d���e�F�������*�k���]��(���u2���� ie��7�p��E�|"��f����J�ka=�`h����n�d{5ҋ)�C��4Ϳyv���oo�gP!U콆��09��u�F�������aH]E�ƽ��tlOy���jeu���R.�����#���(fjx.�7:x������Ä��:�e�/Z2-L�j	v=�3sV�7�q�V��S�+P��J�Z�{`�+�0,����1�.u5v��.v?�gpw�!��2�\� ��):��W�ލ����*׷ԩ�b#U�X�za��;r�M� �ΙhW'�D��	����U ��c�^��{��Եչ�����oˑ�crE���7�L%m��A�o�B18��N	7L�O��%���z�1��9�<G*���7�����uɒ���Ē�v�����}��f/`d
��
�qu�V@f�����r��zKU������|�!0}�� ��+�����/ #T1Mh
��ъ��y9A���u�dǢD6G$'�D	@x��K'��K"�h`li�M���E^�PV��p�O��.z���ކ�A��$���֞o1&�8@����G�9x8I<�(�(�]�=��3yC
�&!�I'�5�mEi��\�����.`)�5�/ocUz���ɸA�.�)9yA���j�`�"�����X6��8��,�)�pr��V�-t���˶)#���������)4!}����Z�n�� �c,Wc}��`t�
WG�#,V�7����� I��_��zԧ1��C[��P 9� �A�M��y�Ll�I�~���ܾ��x�{/]�k@��t��_<��)�����T9rm�y?ZҞ?ʖS��xϑYr���/�x)����\IZ�c߄�cB�tڶ<bCG�h^�*]��|T�^O��;��0�.T��Sè]:�"�/*qHMf�m���X=^¨'ު�u߰��Le�$fZ���(�Zu�h�i��y�Ț��F�3mwru�������h�>�CkZX�g����M}Y�e���qwꐪ�K�+9�Pc�պ�`���U�.�t$�1�i��t,+7��LX.ۆ}h�̐t=������'CK$���{����Ff�kBpǹ��$���)����1��Rf��I�w�C�����y�E��P����#l]5�t����ZL��xgȴ�E�|���!uީ'#l��r�k������wS�Ek�������B��1�R�Hg�$%0 ����4��p%*㫠�F�љ? |�������0梵k��d�c�y��/�
{(iJJ,�U��C�$9��v�И�3�r���M8�yMMN�ʓ`��f��3�xߵ&�j�N�8Nu��JZ��Y��3�kT���B�=��;QSW�U����i8���W��8T���׺�1^�t�M��֟A:^��F��^Xby1���"Yd��<�;��v�é)}�/���L�yy��!̀���۬Τ��Ȗ�!��+#�Y�JSXk�1�cn.B��(�ʮˠ�蚭��8('3�1���V�_��
�c�Gb�HW�c2CX��^»��
T��L  ֕|�l��+��9"�찧}h�����w+BA �"��ṂB/�&
 ڣ���Fʁ�o�9�B���O��R�ŝa?�@�X�DO(�a�{*x�V)�� �̪���E`��X�]4�)CZ�U߇U[�q7I
��K��@ �3M��;�a^"W�z�� �f�s����PM����K�I(#�	���1���n�j+;-�����A����~_���������b���ަ��i����8(;s��&L+���_9����1�Ukm��[@8Kn��(ܡ�M&��;;���Ca'OC��4�����ը�r�6��/��-�刳�u��^z
��4�/3�|����f��U#8Ƙ|:m�� �_�z�x/�/�n7K&��8K�
���p��=�j�"G\3��h��$f�?��ò����׿�d��Kb��wZ���������ٽ%~���)��!R�C���ؓ=���`i�f��L��TO+�}$��1d)k�3k֫m!|��=^u��:B��l��6.P�+MO���Mu��#�e;���$�s))l�ǂ1�<3M�n�9�|B|�v�2�hv	����`������'���Cs{	����F"5ծ�7���Dt%o����dO���}��d_ʿ�Pb[�59�h"����8��1`aQKJHDb����o<����aP/�4&�O���
RBg�O�s�b�C�ȧ���П��0�ׂFӽPO<�����c.+,~"�#u��uX4��)^�E9L�Q�Cf�̊�h���g{:qD�����ܝ;��n^�~�UpC��A>�"���UBՒ�����<P]�|��}fZ_aܾ�Ag!���o�+ͱ�|ȉͭ�vt.���g�{Ɍ��B<���� $߹����V�&"�Jd;����H��󪆃b�h��F|S�?=�S}�jv��� ���*9b�m�I�E�K�g�U{���Ѐ���z�4i�R��iQL����'7I.^��+�	f�V�r$�l��Gw�Ȅ��P�����*`����3j������W��_�� �o+��h�9���T|�b]ׄ�0���7�$/�9O�B�(kd-�e+�bai"U�E���Tu����.��AA�ô0u3GB���T�hC-���C:����<%R \���>����6��qv偱�̄�z�ח,���L�i��H��WO�ΖR�\�WI���%d����u1[S۬�/鎷�r�����$¤F(쭍&�'��ؘ-�Y�}�� Ю�ǀZ+jT�,�c[(�s���˸p�l�@F� �yǱ~��k'V�{�I�9Xu���W�.�*����|�X�b�)~i ���I̞�V�;��=.P�����ǌ��ЬqJ����N���0Y-�pW�A�,:V�� ��vg>)�B���8�ź����JCM?�������?!N�3�.H]>��FL�N$`���M�)k��R�:��%X"�[�Kk %;�JX�~�뷐*���c�?�6O���׎H�jN�A L>��𴂰��б��4gJ	�'j�J��z�"3`��KL�H����w��<���)`f�N >E]���>�n�N��:�zWV<)��)e��E�J�u��{������$$�pOtk��%��A����+W~$����C���b��kY3I'��Y��	Gk�~���h���D�mBjݝ������6���6/m�& /���G����Wb�?��3��g���|m�]��1�AϜ�i��n����ME��MY%/�RI�l+���N��a�e4�lu:P W[?�߱�Tƣ����|�]��UY����cԞ�uu�7ܖ	g�������
[�ەV��`�[�b��n���'�d���M������Ѭd�(��i��y"IPfJ)H�V!�;梌!��!��嚥���N���� �:	�(/.�"pԑl{(�Y�
,4��c�=
ȇ=� krS��*�J7�(�֝d�Y����L#2<ᓗSoe��m5���KUm�[8� ���	U�TU:�ѷ��˒�TB5&��qg\_�����
�N|J�ӭDy�ڲ�s�i��P{��:Y��q����ӭ���B���!��BYJ�u,���
r,��[��9�9�KE��CR*��V�n�;'���y(��Q��9v9_4������C�c>���n� �0
�ue4)�(��8�f�-\��C� E��h~���m��0��m/z�8�;͂������F?��M�Ӷ���WI�Äcq�zn��7�ٚ8�E(�=�bK�Σ���������J,vE�C�J�9��q����7pQ�'��\n�W#�L{�I�4ec1�x|:k+t�	���[���֑70*����p�	?D%%��N������¶v+�V $�$:���޼���*��4]M����Q(6��-d��l� 	y��Ţ?&��٪{p����" �Fs��	��T�rK�aR[+e�҄�,���薵H��BPT��cSL�:EJ	���J��\C�m��1P��,��d]�y�"�I������騨�'(6��b��/��X�b{_8�O����ch�[�W���8�ذS���aܟ���+1Ϯ~����5���]�ʙ�;��[bCV�i9&��4!P� ��f6S��	tkaM����2�bh�"��C�4D���__�1�=�;-q�k�1���T�	v�!B���v�)����&����ȇ�����@�Ź�r�A4B"7��P��@Qu:�Pw����`����S5b�۩~�!m<���F���?$�P_�e�����(	�s��X�Ɩ`���ā��4?lf��˓��`��l��v���q�Y�N�gBq1�������Я�S�K�����jdo�-%���g� ���!�F��{��»h^ҭ��:�������hA�(��ki_��uM?_��7�$ܗa#S�W#⨥R�'͵gܹi�dx�!d��z�L`��ryhbL)�>te4�$5[�L�8`����s����*m���%-�v�e÷��!Y�յ��fb�;��� ����~a��wĽ�`�,4廠��,�ur�)k6������� �fT%��c�7�����j�3� ���rm�!��u�?]��Չ-��L�AL�$j�oCC�Ht�&*/�����*�H�p��X�4.x{��댹�y��hU�)Ԡ.��Ι�2���K�Bx�d�*��h�@�'R�� ���k�~BҊ�g�hg�YR�}DRm3�,�I�_~�m���U���}���W<2ء�$ZcÞ�����X��<��y�ʲ���z�i�Ù��-�qj�����oM)�蔴��C�6��牥J3�ǧC�c]]��ЩH�R3� �!�8I�J|�p y����F�gcp0�ˬ�r+Y���s��vw:E��V��]IG���դ)�q�������]��
���t���3�'E��g����~=]Yf�B��ş�j/�)ݼTe�$�D��EL>L�������I��~I��ݾ$��q*��m��H/��V22[��]��"��g�.�������dE^4�h�I��hC)�0�ʉ���ɤ�%U����Ķ��3��]I�S��>$)e����[y�Ϟٲ@�Pw�z����/�e�_ԯ|(
fȿl�0/���9�&Y[�\u��H�����er�4����9�q�f���XG��c	�[0{�~���I��?��y7��@b�G��q)ڜ�ҧ-X��sR}�[���p�I��n�L�6! @�f	����R�G�.�='Z���	��O5f����쿥A��z��I��8�֯u��X2	4�1	�b}�}ݎ����F�&r{��u�:��Ն:^,��M|j��֤�c�LrYJۓĂ.w:ǵ �8���tn���!�u_�h���YN $p�W�}"�"��۬�X3Êө��d=���GG���'��G. �*�LU�8�e��;��~K�T��H��>GY��[��e*I�~u5~����:�����|����&����z%mm������ �_��I�&��l\��x[���]�h'��Dt_���a�H]�e��s.?�?�à.=�~�1I�^�ʝ6Β)T�L[���c+~F%Ռ��V.LI�H2�iS�Ī�V�Z\����b�*��;�
J��KX��U�ob�s���ι��Ls��\��Γ>�o\���4�T{��'�Q���� ����c��B�ŀ�$6��p��]���v2%����S�1���Yf��I�MM��Ӳ3�K}���2���w�|��Cl\�v)�+��@>��5��Nqx�k�1����)�{M�ږ�!ɿ<�s�,����W����j^�In��(.`+Т��BF`g�Ѓ�!���b:�Wm�b�&��K��S��N���_�]Ұ;���>˒H`=�5w�����BIǎ�ı�UҨ��6\�������w�P2T�#��=�E�3CZJ����kP���bwu�#zXySIjHo�锌w9>��U��>K9S�%fi#3�<�pcɦ�8�	��(8��̃���4���20FD���,���4��\�fj&�b�R���ź��8��\�� dxB>01
�+ߌ)�產�:}S��Ŀ���2bI�3'2���$�aD���16�a	��9�:;q~��4�vӉ��@���0�೤^܄�����DщXY��U�^B�����L:y���X�Evi����ȫ��fL�+���b�UA��̑7�i�G���YV�L�ҥ�=�w^��!W�썥����E�ٲ'<�g��Hi�ˡ�P�/��Q��0�21��6�����֣!����ڨ�yqU�P���M	�q.d�����͉F�J���b��yU��cB
��K�di�R�Y���ۢ7�}.f��

�h�C�iKq�0'��l�!�QU[׶٣0/��S!�Dn繗�����4r��?-���Õ��-CS���Y5��Xi�U.P�9�y�_��#׽)ZŖ���gV�V!�0��6% ��i�t��TC\��zE�ǜ���Q"��e�������-�5�K��h��ǣ0r�)-���N�<��|��S�3�p�_[��Va�7^Q!�������i��y�/�{�Y;�	�X�w��=x�#�6�_�D�(E���T+!����2�Xr�\�䩮����p�Т���i���� b��5go�3��{�~g5V͛m���iVѕp�G&�$�@��2��'���F9OB�2��~S�0ѽ)�ŵ�Q3qV3B*z9�!�X�*{T_矃��b��P�7�������K�Nx�"�rO�'3�n�^DQ�Nw�����ѣ�4������e��zZTA�����X+?����8�m�Qt<#jLeHڲH6]
��W��Aw��
�-�W	�qR�	�"�������K�_^��ݎ��0P��S?	A4������z���G�֦�6��pba�&�}m��
S�wp����X�4�s���9�b�2]7W`�D"Ӝh���ܝc~pD@8�k}�L�ҥ��+��BڜL/hM@)7U)`��䣄����EF(/D#>Ȟ��	�:�F�����X�Ɔ���%cG��ÖF5�794&w�n�ŝy��
�ѝ�QW�<z�Fd�	��G��.0&���gѩ��TK�e��\���K���Ц�)�dL�=�P~m�3�RÜ�CJ�"���mf2#=�����d_[�S �s��-<���՝_6��b����s�@@��������s^�b����Hgu�����˃6T4Hvgz��{�h��(�ҋFd��OcR�����|��)��*�mmc�!52>s$sGb�VUp��4�Am΂v]��_ܛ�p�]�+���WI��Y`A%Ü�Y�,���'1�G���?�x-z.����G�K%U�;N^��Ȭ�="��N��f��'Y�$��i���6w��	���u��2�}�&��kcE��7!�3)�Q��s� �K�!E�M�[ɂ-�u����H<R��~U���WK"�{n`"Y-G�����ɨ��hWB>ZF%���=�w)�MNa9��D}�2ƾ�h/y�;�1�|���~�������s�b�%���N�	fF�� �I��S�o9^�K�'�5�py��r%�cƞ��z��DZ8�1=6�>ۮ	�쬺�M�J;��lV�htRf}/�nKE��8;׳��d���fJ���]�m'�1����C���ck_���q���d�#�S����0`�r�E�.���xX���)�Xe�D���h="�L�\�����q��!�e�5�=-¥hx!�lW�[�sA��٠M�]MB�׫U��j��ı��,Q��k�E�)4�;a���2�7f��)Md�\+���4���}�'s��Ϧ�m2��u��`������� �,�-���7pq�*=s0,�M����wBA��KV~��L��Jx�<Rt=�.����LN��G9�D��'��z��`'!�j|�+���9�<�����{9y;s�Kΰ�9�b��;8z?�e*<��4�﯆���͜�S�qT�O]�Cki^";?��͛r��#C?�=��x�i>M�])1���?��3s��J�)�}��1�q���

9lGL �:���cp���Y���(��O�:9�&ph>�@m�ӆ��@qO��!*3�QS�� �I��w�o�� B�]�+eӦ*�1r,� V�$��W��pX���S�q�4�pY�P�|�����t�����N\zI(��_��O&5���a�q�7n�,���cT'��Tg�*�<�,� �l˫���R����_Њ�my�k�W� �զ%��?pϹ��=��U�J�o��=S�o&s�`{��DWYr!�6��ݚ�z��.��%M���R/0Iڌ��`X�J�V$l�5���}���p�?]�rA�|T��p8Vt�e�H�4�W�u�&�1�UF1r��3wt�ֆ��S����7|�x��r�΢Hh�I_,�}5�\?�^�3���E�!�z�B�@�0�R'��C�(b��3l�'ln�]e�I�X,���]���e�GI"$�0d�{�aN/�3�+�'x�|?�w`	3��8��P:�C�z�����J���ek��W"&W��%��E6�9���*�K,�R�7I��$�j�/9�#2�/��Er�x�fy��������D���H)�\�Z��H�������<�e]7@�h��O�"8<��TI=Y84#�^�n/��:�̺�u͉	������[tM@bϮw��J���n��F������.�Do��ܯS��55�3F�#�=�Ci�f�(W\�>��(��RH)BH�/�*�4��:K�����t��-�}	�ȵ��nz��Í�C� �p�0
��0�徳�IA���w�P0���_B70�چ?�wX������J��Zc{p�K�sF�B&9�#9������=GP>,;V���i͑�m���X�u
��, ���Ի�J�NA�V���k�A8� D)
8B����ͣS0פ+��5��������?������1'F�eA�`�#������lYd_hݰ͆14c)^T��Z��6�l��*�ͷܟG�L�������!���3嘩�	n����u$a���$M����h�c���j��*���Y���!�t��`�D�8^�z)N\A�O-�H�Oq��ŶU�wK�\�#�0W� q��'n�co�!�S����(}5���,zV�+�F�7ҟ�ǧ'w�.x�L�g��h���F.�X�=s�l�^�}��&�=�.��mꪑ����7<���EÑ��~x����B���9�6b����<
�r(e��A��T<B����au-�;-wZ��ש�w�E�n �O�$i����`.;�6ghZh���]!�zT���Y,0�Y"��jVAc}�x=%�-��*l/��ψZ�5�/|i2D���,w5�ˉ�jX�]/�j+n#��\��"�{8�������(�"����$*jn�M�x�S�mD���F����U(QUR�u���$D��T�8��7c�A$��d�:IO�>�(*MY�f���3k�6� #��F2a�c2�{��}X4�W�T�[*��,5⇂{;+�+Ql�#*�H���)�V}�)��/��G&�%9�MY�d��L	[��b˒XMmB�����қ[7�8�,���/T�5���"�%|��ݤ��y*�p�DQ�6piVz#�����=�p=v�Yag�ۣ|nU1Ԋq�4�2s�]W��wi+.@!�L�",C�l������EP�D�������Ǐ�T��Q�Lr�wM���]SZ��&XybMͻ�?c )�J~�Ȯ���bq�C��2�]$�YU�]��!n.9���_ǩ=�Dy�h����.�tu�Y��mbV��`���T
LҢ<S��1��X��,�+W���5F�^16w�A�=>p4�J���߇�(�Y#,�~;KJZ�ޑ��|t^.�sU�>���"����cu�s�yLzŚ��O�:$r�qq_�Ip����"Z����|���v��?��j5�,�#����\��Yqo�_<z�7����.Ԇyy�Z�m�C9�m��u�O����?�8��s��2hH�Yp��#ĺ�_�? ���L���M�aA&�8��#lڵ�,>q[�
���?I�1s���@� W�f(M��NM(W	��z�m�rf�`�V��z�c�r��ʤƽ�]��dR?�R�u?�	�
��~���r~���c�Ke?��~$�8�:����dBE�g5���hgd,ޞ�i�֒L�L.E|�l����,�/����y�� ����t�\7qN�?\b&}��6��߸g��k�*
.1�
f�_Ԓ�r�����)(���|%���({��л��a$b��c�X܅C�@	T�ӆ2[��W�
8��Z-λ�����k&�TB�����P/A���w7�Fd����f��X4t@��Fj#q���ުp(����zBF��~T���#�F0j1���.uo��������B���4?�R)G SP��@�N�|X=�Q���s��|%�R���^�ΰ�@��	t��9(P�GU%3�:���!_}�3m6N�a��S����ђ�:����(:��;��YYP�o%�(�%B��e|a=���Z�ąe;����~���^*��6{���v*ҵ������m�꽚>('*�YW�N�){��;��>^C}`QV��} ���iWNe9��'�$�f����Cȷ:��דf��^�Ut�! �L�ȫ�-��t~����fZNO�7BG��Ξ'~�'g�-�'�jqL'a�kp��mK[�V�z�]A�1���垕ſ��c��S�'!���B�_�����h*�E�b?��Qi?���!"�,�-h. Jet?��=�5'�t���@z���D��Sϼ�u�K]'�ď_���v�O�����P!gi�l�q�Y��Z�Y�b�^E��i���W]�~�q�L��*ӀR��3��>�5�z�e�
��S��7�@��?�����0�j�`���
��i���|��$����;��y�|�Wp���(]�(kҺWv��R��y�������y�ᛓ��^1q�7)��BRΰ��K>�|�����1��:WC�a�>����H�ɇ�1���^��l�v�_c�p�bD�2�ۡ�v'\6�e�/���|ʏ}6�+N�~�ⴋ���~�e�qR����:w���p��?+r��o��v���4�wf�~��\̽��Z�:�Aҝ�-�
�*�����
5#i�M��K�~b꥕�v稺X`
�Hr��oX*�s��2���֓���>��%5{�m� N��*�2��O{C j� �j>Ȭ�e��>��g*7�	�v.$��ZS�!a��Y�/�
�V,�L��[�M��D�=�R��{��a��H%;�]�F�h�Q��`�����h��z����S���7҄�g�����[Fg���ng��2ZŬNIO�$g��������#A���#�ǁ����&o|��w��=��l�'rY��ٲ�@���ؙ [{��Y�,x/��
�ě~�/���o܀� �!�lH�B�� ����Zu\��Fi;�ߠ>`�����`+u�*� ����T|�_�V��|�lw�|V�"y�%ͧ?N*rƸ���hvd��8"t�	o��~̹>"Rn���Qf�G\��,�B��c��!8Z7�o'o�D�B�d��R��0=���f���ݙ�V�\�վG=�{I�i�O9�*i�C��E[$Z_���mc��B����압r��H��o^���k�;aٌL��(?��Լ<�z����
��̐��o$��8�38:�E��~��1I���YAN�&E��Ne
_�i��k*z�V�q#
���5"l��;��7�w���4�c_���9;�LJQQ�T�e�m`]��X���L6��H�2�;%���I��^NJE�N��	�;c,9��wn��6Ô[V5����;�f�lʻຫa�U�Q����e��%Q��*-~˞c�ѥ�V�%G1�M�� :�p^J����O?��S+��Y1�hC�d��n׷?��-��RT6��R����9�n\��y]���84D�����uF�@�%��9��#��C�[��1y/�X[6����s�\�.�'�����>���Z����H��1�����6i���ۈ{�$Av7l�u~�.��W����5��}�����+~#��]g%�t鵱�0�s1�t-��9��5I�5�h9�%_(��0�L�����DeD�S'	g��m(�Ż���Ė�n�;��ꦺ2�8��m��������K�4����yDՁ	��)(t��<�5�q�nDQ;@70|�M��ll:�!�>�w�d������$�l��iT��ݳ
�0%�������z�����z��͹!1 e@����10ds��#���rS�z��+&*Z�C��vP��|8��W��1i$(Qq��f֮���h�y� ,��qL����8�Ս��]���H�G�UGdDe9p6��^C��,Y���*�����Ӣ!�L���Z�^�-�Y@7��y�Q�ͨm����0Lr?�t<M����z�!��$T���F�u��Q8{f ����8�����4��عc������+!�C	b<]��ô�,�b0����ܖP���ơ������JW��b�M�&"�����w��xi�Q�S��a�*�������h��u`�S�ϖh� ��g�����j'�g�3H���t����c=�aV7I����]�������Q���ς�b��M��&��5�Ș��h|��I�����=�6��͝f���ʚs,��4E]��zN�'���ʮ�I6'�mi�Dy�^:n��h쾸%������i:�+�`��|i�Ak0a�C�;�����+���8��$lxU�Q��T��H�9��&;۞�mS��_9Jh��zM.6���o1x"�"e�T&@|4''��]��|�>ˌ�9Kb��#��Fk��������ni3���|3��`F�~�ZF	�'ˢN#}8�6U��P�&مbO��c��~B�;������A��ΑK A�����~�{�O�?�ޖdf�v'����:�ٻSh�R�W�߶�V�(���Fj�B:ҝb���k�c��2���lXX�Ď�}��M ���>�f?��i��v�r�`=�S��ߒM��{��8h��
2�#><}W%�s�_2 ʼ� 6� ����3+$����C(�J��(�"�u~�͹�^��5�A87�:XK��}D �@�9�˲�o\+�W��^��3L��z�*D3B��8��0�ϙ����*,to�TY{C)b�v�[��LǊЫ܀)�x�V�Cֺ�I題��mG8� ,�^~�v5���ҷ9=�j�s��4"��|����-R`�M����n�c�u�M���L��i3�o�)�%�Z�����zے)���UC�ZL�$��ª
6��R횒�������c^�,~a8Z�]�����c8O[��e�c�e]X�1Ѻ�/���'hPײ�=W��39v�����h߉Ѡ�Ȳ�n�>ޖ�-B�N+n�!��R�*]�#�II+�~��xn��F��;�ź����Hju����
(��{I0nb�� ��ھrK��o�jJ$������s�d���"����9xv��IAf��lVZ����Q(��	*B+���-d.��d85b3� E�k�Y�ӸUB|��j@o��a�L1�S��CG��ꆴj�R27;6�/���}�c�0�
�R%֍2BF B�ת�f�!4>L������Tס�)��������mg�'u�i|oV�Ә��pӟ�֡˰����QV��05�����Ӧyz1N݄�SM��:r�$~����@�k����Ј^۰� �w�������-�hZ�m����t%Z�Yi*�t���!����T���\־�p���-F���B��Mع�_8ibH�Y>P�[J�}�X�u�ʚ� s�����)���V׎�Lq��� z�����d\X�`6RQ틙x�zpZ���m#b�ɘhⶊS�D������"�4�<���_�*TwW����S$13�i�EY���D��nH4���A�S�z���0%Ƌ6\B��������fk�������M�J���Ȥ�1�63)i�ʶl�`LY��n�\��{H�����=�)���<�c��Ƭ|�`_�����@���	�"]��8�����k�e�Lo���1+ΗL����D��g�9�k���lt5�e�n�vg�̗���S�P�EJ��m��d)�9G��K�N:-�=� �t9��.��k�a����?G�:ޅ��L&��]�wm?�2�������|�\
�X��(¼�	E~���&���J�\$齨�:�n��a�,�*-����;� lm?@��~�/lٛ�ݚRU�1n<4��f#�|N����'��	�	k��a�y3��$pĩ���
�/QF��e?:�G��i)ڗ�m��&�q��}��g�-��˜O����u����n~B��C���ŕq%L\�q�|�������N���Z=CR�DZ��F����H�t��;�2��#�"
R"t
΍C4�����q@n��2��5���붯4��qZka�'����>�M+m��y���,DN
7zk�cy�I
S����7(���i��Y*ј9�	EJ��nڀ��u�A�=�S�z`{%����n�Dn��te�^�xxU�<�3�}�%��ȋ��0�y��f���f�kg��o�j�4��Fi++����H�֓�h�#�u&��n"w��鴖"�o��'{������bO�*ew8Ȫ0l�m���87�1d�������@n�P=�\���K1DG�mb� D�9r��E�d'z���>��{�:�0���XbW̦ꋊ?= ��ʾ����C�K�f,«�X���K*d�n4�KGj̻���������熮�O�[�\_�}I+�,�LwJ�,�ތ�����곯awr��e�LJ�}�ɉ�$,��N�o$��c�T/��Dm��s�۪'MO�֍r�	TʏL���8,�������G��!�}.�ۘ$4U� �ԇ��{_g֡"�~ ���o�:k��v�K���Mb`V7�
���AA����`�H�R�'1m��O�nJ� ��+)�`��V���W���eT�#��l����|�3�~4Ƿ��[��� ��%.��`�NQY��R�4+��]��S�F�|~��0|-�����aնȫ��'�|�4�%��B/�#�<i\��g���p�]����xq�+@ԟ�W/���$-���b�����lb��H^���}���� ��(q���yt�Ⱦ�+[!B�aݩ��a�:��uY:4'�~Ŝ#��bv��C�4�Y6�5�AG+����`�R�j�?m���[J��B���/X��cq+a�l��{I���'��u�A-*��.\��|�(��6�+Y�e��^O�f�)ҷ�yp���f����Nؘ?%ʮ�A!��K�j���<&��5W�� ��t�niu��U�Y}k�i�E繘AGF|��Z#'�2�Ţb!���~�G��F�z-N �3����
y��$:K*9z7��B�u��meY�^������_��P>Z�VN
�O-'���V�o���_i+�7��-Ͱ6T#���d��|ӻ�>����# �T�C��O�[�'W�ɧ# Q@�T��� [�_�E�?"
��4�6��?��|�#���q��C����8I<}%���f�I�Y�#)k�'0ؕs�A��?>�1Prx�팋>]�'
�8܇d�`�аx �m�L���7�n�/K�ʴ ˱r�/(ս1�^6�x7x-�);ո�kBhq2�-d?����@�yLx~�6=yN�8�f|U��c���#�<�[�d��#�H� ��Z�p=��*��&Y��:y
�<.�D�(~Ƞ���.�e��+0 ����nǃi�~�"a��fQ���W��-?v��m���S�v?n6���M��>�7��ܒ�pl���^џ��.$��\ }�����%���/ލ8Q?���2+�*�g���
ҡE#�fe�g��:�����#�?7J�&��q�l�|R#�>���'P��,��X4��X�y�uQ�*��?%�,R?�'P��n}y��%�f����Rm�w�Z�>$�������j�#����T���6?I�[Jt$T��觌V1Uq�Cl%�.���u*eЀ:><=BG�eL�i�Asݥ�*_!e`[���)�d��d����q &�Fk"��tr���?���P��PR,4MI��'̙O6�<G�*���(�B7)�<c��ɞQvL*�МQ&\d��zb��M��|DC�U�P�ټ�9�m֑� ��%YpR�}lZ�a���#�U�������i:9݉z�HVr� ��<0�&��$��4�:O�|u�ݽ�7���"W��5����:+�З�&o_�Y�)Z B2M˂E ��.�����rŽzá�,�Mt��C�$��{9��@2A�M~2��"�~&�#r��'o��2?���b7�I���L�#� �c���r�2��F�'�4ut� zYeQ�N���{��f}�OA���~�G��U��~ ۥS�D~��U��>4 �5XG%�+�+��'Ь���j�I@���ԁ���:"��/�UMC�0 p
tQ�`��Lsj[�#�C$��18|x�z��*'EKIK��"�o��qK7P�� �����6gê\���[i?6����znnB����3hE�HX�!��Ȋ���.=�7��Hh�5=gu��(�����A�mq�m"��ݓ��������F�;�S�;q#tm�2?`���.\��
��$�j�북�gr�]����:	U�⃧�;�!�ZW���2��!83�8�&���u�x]>V>)�^�i��&ai3H����|� );���G�j��HEuTNkJCUN��|Hj���:d�_�l������2��U�35Eu
vqOY���cT�ќ��Lzme"ʈ�f�yW%:�"</F�YU��^c)ⴎ)���PJ1G�����H���}���\ѻ�U"R6�!áI�U5�T�K���� y���pEO�� ������Ϳ���N�v&-�z�3{�� Kl��oߍUڠz��F�;�=%���dƭ�/$�����p���c&Q��ϥ�B��� �i������e�}-47�tH91$��$]���V2`ڴ�<ӵ��PV�xߩ�:�[+oM�>W��sm!�K`O8��FE�r���F��Cbǵ�^�aZ�������;��Ҽ+���>���������L��E�[�����Uv�FL���̼_�J����I4�`ҧ�n���ӴxN����H�x���y{U��ΐ;g-ޗJ��N�x�Ǻ�՜t�`�|�.3���Z��4L�t?�G�����}5q䎴$ꪓ�¶�M���yO�8�\�j�����!_��m�+�9�����p����9#S'�KW�ʹ��1{�Tf�V�P����x�����o�{q�|T��P�ѿ6�iuV�s��Ї���
�㷸��Pw�Y[j��s����wd��w;��׽?
�h�1��.��䟃��$���V���z��(�`6�B��/�ڶ�M*�'�c��F�oVj~M�<�+8�!��]/! ��J^�|
WC�x��i���V&!����VJ�MF7A�wy�4�p�����lS%2�a#��l���ܛ���8�,A�:����n��`�2.}2��%��$�}#��/��X1�m]K)RV�.�a���?W�.c�|��j)�o3Q� =���Q�3��$P+�0]�pQ�:�[I����Ո�UTw6c�����ϐ8$a�d�G<�6��%�\+êkY��(�d�T��	g��p|Y���fOv����E&�	�sX��C���߳K"ް��K��EڰAh��uȺP�}8We�$��(�G+`,�v�57$��hb��k:'���+~5geL$nD!.��ک!��͉��0�^���ʶE��~��h�*&�mcK&{�6�Z2^_����y�� oB����	�O�,@�����~�s](���%|�k�<=��.��T�����Wk~��IF��w��b�w��e����vg�ϸO[�OE���am�-&����V�����֠����sJ"�ń��E���Ǒ6��5:��6|8j�<̀�@ {�@Z"g�<�4�k9����6N3BU�a�D5�=qq��v��$̲^\�~a_�d���Z_��S�!x�(����׈o/56�&���ó.7%c-�5�i�DP�Q���Z�x_ܧ�έ�k������|�;ea��A�O�C���(�\1��n�z�]Ȓ���tU�~�6�+m�s�I=���+�)4�b|�G>1��uD-b�j0�G (��/���z�]Ն������q¿r;Qj������7~l��V��G����(ƕy�����
Q�i�&��Ы�Y�
9�<��N�ȩ�w�ʘ�uyb��Q�?�HR�M[����m�H"�U^&���m�����"-��?5J�r ��ɓ�֩�8���d��i�PJ ��=�y��o=a��L��V40wI�p{����,�-��f/Z��=�{���Ih?Z��e���sH3>*�䴋��e�k��P,��*����Hχl�}�ܨ��t�7]j��˻!��6&�+p�fer��j�h����<�Jk�4���*��^�3c��)6O��pn���c���)���T��~���[�;}��EMۦ�7E��=C�<ur����H�� N,\�d�¬��"���0f��+�{��/p��D`}��i/?�Φ��w�A�h$3/�Y�L@6D� �i$�Qg="�r=�Gۿ�k�r�D�l�f�{�����޴ �S��Gd?_�o�J�<e��┱��p2���s=���b��(-�
�9�ew���>���?����3Z1p��|��G���P�L��t�.C]N�Ʋ�0���p��t�/���Tq~�������c���SqM�$��w��t;�Un���'�X;��G���l�Uz�1p[%��B��&V6Yx-����)t��{㲔G�y귰FJ����l�O��rS���W9W��t'����z�&�ʧ�T���@s"�VU�	������%���Z�~A�T#sƾ7�r:�����iQ�.Tg@��b4M��/e��|�csΠ�Hc�I<��p�xJq�f�: ��L~D
���z>��>8J��_��<�wlY�]� �Ңw����3v�����tWwl~�� _�o��!�o;���ot�,U����9��$�<.� 	�.<�F�=�'a��s���4q�����{K�ީ`b���K �1��]v���~8=j��"KAwb�8x	\�]�$����7#f a[���ᙵL���9Ef��Z���z��S2|qHh�~��#�7�f�T���(�Ӊ�^K�Z-��{��VşJ�ʪ�6��9�Nx����f�V���H�3"3��CKe����aΞ�{��Ww�КI�VJ?�&���R)�f� /�B�$H�2�Er�B^j�`ߣj�1YY`c�?��:E+R�ӆ���=��l�B%�"$���kaHʽ�Y�q��]w����wa�N�o��۹ +�]eG��_��S��ܔ'��e��;�����P����[:c96��E4ޗ[E#�2)P,��wq�~d��G��A�Z D�>���x��h*L]l�?��7�-����b�Uy�h�����k�|jN&GP3ΚQ��(E��AM�w��xb���)�_~uW;�j��*�����rA���d�`������^A�y����
B�c6x'H�.������R�%�B4aG��7�"�Xل����,.��Шćw�]"�q��3>�� D"��K"L����l�5u�j&Z\�k@ٺ�+�
�T�.�u�zط?8�;�6e&rZ^;O��P|�M�JH'�gK=ݯ��r$~,�C283)|(�永���pu�c�=Tl.��]������c���}kb��VF��|r��+���$%�<� B:c���[��w�V]!ɂ����C�[�՜�5S�4��mh�r
3JA�Җ�-�P�-ڶ�%!M��r�pq��6�N#�w�<	.@�
&�gO�w����ՙ�`Mhڼ��˫�q�E���J�d:c0�ik���W��l�"*K�Ю��
ٸ�7X��-��T�������v��IL�Ύ,5'�roɸե�%�yw��
l��:�cz��J�����$�^�x��� ���{���� :�a�P�
�m���&1�Ϭ�[���6	l�+������6!+�5g�ͥG�^�E�+�憐�����옩u��r�>�v��|~ܬݯc =�QVc��d�&��S��Q����\�@���\T�ip|V���&�X�W۬M�O[j`8�������N�]8��@Lh���,�*J��2A�'P�r����s�I�d��g`]�ҲS�m���Kr8Vd,x�Z�����l�H��o�.�}Y�uM�N���0��r�y�s����k���6�G��U�A�S��`-fw{i�Z:�����GMu�P�V0��\c����#D׳����@�2�Cu�7]�lp���S��gO�N�A�??oE{ɗ���Tt@uW~M9�A�]{Zz��&sY��y\���@��4��GI/�d��������GY�yC��x�����}�@�C=λ1�\g���CvY[���8m�ZGDU~6�o\��c;�+�]M��$�<N�L���2	ŲR���<u��E�{~HA	��[�nD�S��f��䎶߹G)p�ɰHt�:�)���;��@�ۙxn�~�z��J{�[V�s_Y3�h?j����t=dq�/�x ��I?�|�AI{1b��%�Ah�p�\>���R�2@ ��1�W�9�Q�^G mݙ/)ث�Y~��[�:�q`��i�TsT�i��r�~Gg�NhR��f�`C�s��ƪ3"���ܯ�.VM���7
���g4����L5��L��P��)<w�a.�g/-���0���+�	�"x�,������~�a3��G,Ss$}�R�z������k�f�q�0�u�����É�Xt}��*���­��EA�f�z{�YD�)�pR+ެ~�M�G ��u�c�]5��:���3������6�9�UL��GRI�u1���?�E^�W���
j0���Z�)���M�?��Ş�By%�R��4��7!i$ 7��d�&�_7�Qdc��-���ޓ�!�*+V����(��� ՝޹TJY��s��`�D�ui����2 E�� ��,dH���˙/��.�NsD��R� �AL�B��r���o&��?�|�['�޽f߶��B�s����W6^ �o?��B�&Q4��#�JLS@�PQs�_A�`�&\"P��5����J|]��rs2܍���m$����;d�a[9��J�Qeb���1N�N���7qiA���F��,�7�8�Vo�E��|cج��X���>�����ig���ۑ�)aÊv�����7-��6�����w@��/׳��+�5��,г�2�P�i7��d��'��xn:Ά�v�{������7��;T����f�����@��V��sJ����5T�ښ��_4Ջfsj��ٰ�L`,�F����vt`�T��x��e'�Q���P�֦��F�h�z�"^P���l�j�nթ7F?�w��*�)RF��%�y�0yjS�O���zqYIo���^�t���4��1�lH	t�á��d?U)'�|�#Ȳ���/�#Gb|j�W�|�)2���q�>s��v�Q����׼���.'
��Px<��y��*��( ���V݊l�ǿ��p"ſ>�XVx��U�7����4��C�S�p��j����v�%�Bh�̋Bs�~cDr�s��O:�ӻ=hj�k�	Z�kmx�t�i~`�B����x����.ԩNΊ"B�kn'���e>�n��)?�\��a����"�,nP��1�ڔ�� l��`ῚmV$�o�d~��=o�ա�U��4<)wgI��ǽ�\?H'��b�_ck���P��*� +ǅy�?n+��W�1_)�l��w�L���H�m�}��5�"Ԗ�(�����q���8H�p���f/��!�<��q�v_b�����nP
�
/�3}��B�����L���)���t�r��ei'�=��sҒv&3�.*�V[W�y�*�o.Z�/\gD~��7b�Y���-�b8ib?�B�wY�*��^<�ǀW��8���6,n��V~�(�vi��%e�㟼zߵww�c��q��@ܥ>��B�Ի�c�k\	G���Vq�7���n���t���U�v7 �7��*9���h����k���9G}:8��>���Xd�Ҩ*�VM�3������7V���� n���f��fe�F:g8IN���)04xx`�NU�f��(��^�]so9\�s�s�˹��s�?�����̈́�����hB�)x!o�a�|A�e�L����[�hn,}_��?Β���z�N��8l�x��xEU���o�%�	��%�� �p2�|Sx6��g%�B�>a�p��}D �k�ɥgS�č�*�d�7�BX��^z��<��ׄ�7H~:ͤO_qn��Q`����`��<�x�y��8������)�����[';�щn��M ?�%ڂTe��ZzC/�"&nx�i�\k��Q�=Ţ+�
��N��<+XȚ;�gI-LĤs}�0�/�ٟ��o=�o�D.h�ͻ����u��y?�Tuc�Y�����d�N�r�� ��X=�|i������_OC��{��Ruk�n+�t�V�ۄ�G>u�_9 y;� L��m9n���K�u�Wu �[¡t��`��Z���ܥ���m�)���\�"G��L��Sx�8G�dJ����v���e!����a�C����T�e�I`Y,&=���) "��q�!�9�8��Nz��7���g�q!�zѹ2�V�H�Z֏5>�R�%+/��C�$�:�'Ozg"��<�qtȖ�� �~��7�l�=E��#bmͩ�G�����\�|��Y��0�Co֙p5�[r��,t���q6WSlJ|%#[�
l?��[`�=y;�2N�A�����M�9�����۽xM�ƞ.H�W�<�����qR�ŭ��v��יo��c�I�0�pGk�i��c�(���hB�\i�U�I���e�O�V!lR�yf�����-�z�n��^4�M����6
�m���b��uþG��
䍰��8����i���I��6��^�[r� �ru�D�����k<n�����2���N��Ȳ���l�f�Q)����t>%<����e��MI��um�"�M��١��T�:��5I�՝��+Fh�`KdsЛ0�b0��;�Øv��<�[����5�tfE���[��2xBi�����\h|�4��Y1^i2i������TǢCI;��*Z�t-V�/A����e��	��k�&A��5��nͥ�����k~��ڵ����_���5��z�.}�1P:F[S�u��#��>S)�D'�P���٫�0���d`9*���P�2��X����Q5���b��m���ʌ�B4��1�`��Y���倈+b谂U��O��u���|A��&|N��M�U�t��2��vb���m�f����J�XSH�hҨk(�.u���_���Fo2)�/A�B�3�0mJ5ի��ⰧCjd~(�S�jrKQݎ�?�Y ��9��%>������բ0~g�6�<`5�Cva���SתD��:�@5'�[��/-Ez��ƚ&�ʓ�s�1Y��hǿ�=��N*&{V�9�0\k�,�
!l�S"��Q�Z�b|�����0�	�I`�����z�F��VQ_c&�)�Ά�d]%=t۫+�b��o�4���+�L���#lqE�U;�c��`��6͐�E3�1�e��a}�"����s�pT�y��68O�|���cf�;��G����w5j2~������:�Gb���������S�Uw��%y*?E��l�E\�t�p��b���<���X���J���0���� lF�I����K����7�i�����5��F��Y��\�V��FwU:�-u�nL3����)�<��Lɇ�A&`p�Ku2)�����N���Q�4>�9�R�6���..4�)<�.�%�/leq��,��FM����w�ػ���iΜ�����UI�#��,�z�{�[_��as�_�I�d�T�u[�mSF�]�;9�'�&��'c��O�F^# ��.(�\w����A�fb6C��3ī����7$�@Q��q�x��.�3Y*�����wo2�"\0?��:ƴl�ݲ��"�"�y�=Nc�n$��V��������^��˗�Gd7D>�'��m��88�׻Ɩ��Vn�^D-�AU�����'_<�vI�b�\�DDLo�6G�S���(��l�$ C��3\ޤKPӵ7�BP.W'����l����\�羚qL�Jf:�"�8��k����ڟ<��P�c�u8L��cB��(�@��J�i6MP5���PfF����x��k$��Ƈm�Ę溢��d��B�"����~C�N�f4�>�w\e�լ|��G3f_�:\�>���+��ֈ�DT�U9��U?�C���mԆ#3�fG1`ִ��Rln�)���' ��Ur'A��A�?ra�	A���5�r�|��9�]�!���[GY���Az���,���w!��=ݰ�+���jf��Z��[1�}c��Q��$� v_�Ä7P-����J���T���B��֗�MD&Q�w�+��fߞ'S
�U;���烥o�7"bT� $��O'W��b��@i�\u_/��r�j�(�j�zi�!]����V&�"��WaLj��3����bc����8�d�e��*]N�>�Gh`RO7H�zW=-Ǭx�t�0�͌��O�3z�u?��W�r|��
 �Fyr�4���[tͷӐ���w��c�5��$�<��1<�>��$1�� �"i�~Ο{x�W�$��T'o �#W�v'�/�(�H~�Bd���	�6-h��h&j@X�&E������Vx fxh�1l�	�4H�Dlh�f���SS�WX��t��m����"�ѯ���L�9ޠа@x>�?�z��E��%g�7:J0��/���ڨ_�_��s���SOl�������/�+�$�r��B�4	[������g)�QR���|v@H��}��62r8���j�p+TS2ϸ��]sP��ӹ�z�i�oP�
�%��J�K��#툀��N�������5<Å��u���[Iu}�|N\����-�F�x�}�%�*���,���*��.�(���w��`�u��8� Nb�G��}�5�qQ!�Ķ�ځ�͞�K��k������y��2_3�ߞ�i6n|�^p_SUY[�)��cn�'��D����},:�\l=�Ͷ��?9���o:���'P(u�k���`��{b�C�E#�u�%��#���v[��=_�����Ї�٬��5����E�(�M�#�ˌ�Z}W{�ۀ�k��. )��M�}񿆻;l�'s%���R�;��4y2O۞8�vJJ?8,p�8KW.R�}��*�k=���q����M��<}7�8�v�+�.Q��3l���Q�E��@~�.ܙ4�~-=�F{Z����q�G�:6�k��ŌO��UD�=�Nk�Ab��:�W�����w����4m�|������*�8@N��
ũ��*���`��!��uj5O�]�}+�H̜�xU��ٚ�oy��J��E^Ws	�Q:ut�bԒ������1�J^��U��H�� ]
�����ؖ� �,fF��CՆ����ۍ9D�ܰb![+�zG�� ���T�ja�``���)O03�LqH��58�T�V��\.���f�>"�\���]{�:��ya'�M`'0Qb�9�����h�M�B�m
��"��4��x�ό���JYE[`���[������2������B���L����H$�̙��}a�vYp�}-��
���D'��F4L�{�.1�b�2G���VQ�����.{�����=���b�������I����e������7���{�x����+�n�%�� ]=������FO7����sG�	2g,cM�h�J5TD@)0+[pPN%�U�<C����0�r(17��x��F���S�9�m�Ʋg��$q��!"���)����?�G������p?�r�cq����0w�ƌOt�(Q������	��\.�Pd�`�7�w)���I��é_a:6K����R�#��{���ClJˬ���qstEN�b�`\a�Zb�HV���*ar�+z��*PYR*?(�h'�����9��$�[�0�b6�=�7t�O�ۼM¼i[���2v�d��Alz�س�[�1���\a�v�o�5��~|]��]�����&$.0���9���T�ڐ~,�L���-�T/�W�e� �����qI9s�*���� z�s���>�Nzx�[Eis��S��������B�I�����T���n��3�@\q�}� �Z�dЙm��@s!?a�[5n�C�3멵!o'�:�LW<�I.,B�B|<|�c@���p:�Y�bL7��-�;�34�r�.����&���it]I&��+	��]eq!�gb3/X�m���b�|�I����z�ڧ	���z��-ޚw�i��y�� q{s�F��8�w+�n�$�����V�T�5&��[�8;�	*@F݃���QES��qR.�>v�6�\�Xb�'�W�qh��os6�m�~�U�RU�F��L%CJ���U,�3�^���]���|���t�!�����G��CSx�1�B�����3lY�:J��Qw���& jrB�����Mp6��<���W��ң�S8��F'��΢�J�H�}���N���[K�6���&�][�eg�o�4�Uq���@��K��˅��h����V�R�k��'�'�4�U��\��(MQ���YoP�-����-��n��
ni3��|���0X&���-|E1�Ov��Q��ْ=Vڃ��F��MHn`|��8�\,>���
c��� q[��Pi>]�C�Q�)�<Z~�ȥc�Cde�)��;��"��l�T"Ioz�z�g��\�G��M���"���/S�VqZ_��HZ�ӿ[<��|Y��R�V�`�ٜ��O:�*��]���eyC7�fUE�дLpY��U�R�}�c5;�̵&-
����@�@q���4) �H�v�h��綊�"���W([���EQX3&���9�ƑR`�w����H��ZVE��{
�Z�����5�q��,�l4̽s�֪Ӫi�,2��v������tRj����I,y�����f���`!�j�iVfJ�?�W�qAN�d��x�������1=W�L��ō��҈w��o���%5��&z�G�}l��p���*��nEt��Y]k�n��pӛ`f��q!/<�[`��&렑XG0�ϯ��~m=&�A�8��se��e���P��Q ca܈S��hU�	��"��-uD�c4�ҿ�y�3�R��=��o���f��'(�'�R�Y!,�ڜy�Ũj��Y����j2f#��g^ �o2�F�j���[բTBy�P3�_���+��u2w����r�=�:�O_욑8U!>��������h#O��y�h���A"c{wÝz��|�{Ȕ�(���'�c*+�d��/%��i� x#}6���$<�Wa|���'���v0��Iz*��V�Q���D[F�׷�E��4,�ğO�N�.����%��o��R@[�����.�-�hm���X(U7Rʄ��0٤_Q�1Z��Y+�&!�UYR��<���+��)��#��hv��1k��y����Tn"�N>����\p�fm=0���$�v?~�S��[i�5Ӕ'��ȉ�=�0���?F\O��)�}��
P�4d�ŭ��."�P��^�s�4�����;lW��[�1�A���B$����~_.S�&��MFXRt)��gu�86�| i�LPg�r��\��&Ų���F�]�����9'>��^5�e�_�� Mn����Y����g�榴��X�z�����Q@׫x�#/U��xyr��,�*G�dD��2�?�Z�
"���\�o��Y����E�b̽�*�^B�љ�U���9�y S���6�+>��6X�}3�h�	��ub�O,	9o�x�V��( >`!��V?� �&��,�1u�ޗ�^�e9ՙ�A�G]�̺�Ͷ�Z��2v�h��Wɱ�k�Z�,Ѽ�[�v2�R�=����%�����r~-�&��n��:Cǫ�yU�}���C�������?��.�MU��w{}Ve!����{-2C��9�`��<�E���1w>^�����	۝;�YrFo\��������ãVD��f䳀�_ecy�d�=P��^���M�7��m3�u�W*��e%�m6M�����jKk�� �M�Đ����2������E'<AR������p�i���9�D�Sп���ڐa�h~����� ��n��������d�{�ΝL�6>&����ҡ�:@\w쏪k�F������:_��l���[v��r��{��O�;\�����.�vн�C!%h4A��y��32-〰���z���]�)������f�GA\WGQU����N��9��0R�0���q�T����a'=j?�q�����8�/*{)�s���S*��e�x����g`�ɅK��W�(�����8o��?>sj]����B�V��{�}qpPS2oO0{I2�`H?༤*a���gP�-Z����B��p^p���QV���Pa�ΡgӺ�g����C̅d(��}�W�wg,'$��O=f����4�ɹ���	�&���]Ýɐ�{Jg��f���# Es��"-�8�� ��[�@ t��N���0=oKhʎ��}G��2z �� ��|ks��&��js�I�`O᧲e�/B���}���~����ٺ�mi�9�Eڰ�6��@�����H���l6퐌�{�u�G8)��Lph��pt��J`J@]�/Lu��)��o#3��l�)�0z�I�d������n)!�x��9�oJ������K�33����8T�p̕�+��\U'���<y�vRF��JA=Y�'H�{}aA�� �x���I����6|5������3o�<���;Ղgm47`{l��a?�������Z�n�H<;���R9��.ƁA"P-�#�~��К�Q�������\I�u��:�b @�i7
�?Z6�w3�B����M��V�=�nE��Z���%^�7�Y�����d��a�_/aD�����"^�������#�g&���w�G�^����9�VJ����m��R�zb~B�vH��8O�P�����W���a�=M�&g���a����>j�c�x3N�:�(<����1�������O�d	�u
M�m�	\�s�G��iA�N�<�5�{{���S씸y�|Iq9��HR�c�8:Q�4ׂ�q�p�e�R�Y�G��� �)y�㚻uNv�d�]�����oOZ��oj9��I���;���)HqJ7���W�|[[/�J0ȯ>�t�W�Q{� mS+��`X�<����E��l����=��y�?C�5v��u�-.u�h�)RI��=�u���=��ִH�M.Kka
�OGn��HvWs��J�/��^U�L����������d��<]��S	S��N�Y}��xy*��	�j����?-����ZZN.�m��3w��}�Ƽ`���\ԐN;a�lz�0��c�0J^P�J����[��6��0�D->�\��"�􀑾��z�ѓ��Y:���>O8�)�֭K�ϐ%��cU ��%�D��o���><�J7��&��4��o�n��T�gm�h��[���[�k���y(׳%�,�����U�Y?W�]�b*?��!��ji��*0�j+��}(�ٽfܣ�c��d�.��\M���w��u�n��'��� �Q���5f�7Q��|s��]r|������l{�,^�RVxI��*I���G6�I�E�c�P�]�{SX#���2�kפ�ձD�)wb� ��hK�~��ë��M�G�=e�dx�5V���4�R�B��.�4vJBC��t�xC:-��5��;+��`^�F�:N��}#�	f�ۿQ�L.�6��CjӒ�u~	�Je�dȐ}D�Iø(����0�<KI��p7
��!�V�Ub�����~�)��|*��r�� V�[���tB:gY��8��O}.�k����j�0����,���&}�%�zFz�*�����o��˱�!�I���*2�y�I�1���P��q�o�;��E��j i�d&�::�4'��Jd1y��{7¹�U3,?�f��ݣiQ��rD��ߚq�����G���v'���ԧ���v ��ѳ�ݍ6�j
�CzOk��������ě����[p�Ǣh�ߙj�ȝ�(�h��N<��.�vp�mGMF^�[ҙ�r��Zr���6�yy�(+��nz�_n,�\�����=�j5Ǖu�k��"煍��V�Wx=xi�類
�!���W�L�}?�(��?x,����:�囒���ܩ]7,WA�M>"(�&G���!��+7���8˩@���P��N]�M{0Th6݈�kft�=�;B��Q���ꆖ#3p�{��0�i��u4��O���>79=9��²
e����yf��O�]����ܻ�6FD���x�h�kj���>��Y[�^��왖4M�h,��2�pl��2;ĭ�����
�?A���L?��.3�>�qք�9=�L�Ð�Ux�+��5�����>H^~J�K�`.>�Ϳ��ۍ���*l�#�M�`�b����zG��Q5Ub+�|���^6�G�n��0
-;*d���_@���*4b8W�*�I?^ӀV��rS0.Y�O���F@��Ƞ�G���z�=�,�[%x��O<~�2],9��9����W�X���I(P�ȬlVQ�7(�P'�#R���8�H- �*$Ŋ���2�Gwý`tk���cȕC���V�ڍv�E�y��,�4[�'�lN�'S$�z�Y�Vf~D�.���-f�e�xn���y�
a8�K�ge3Ad��ե���M$\�Nq�lڶ��ԑ|�5�9�	�^�!�{(J��q��N����0D�L|�I+��sQ�;{�+�6�Pp.��o?Y��h�`���t%�7�>��R���	���D	+X~��w��a�X�m�ێ�ǲ3$ŋ[� �cX7�|/�
xj�?��r]����y��8V�����a���j[ $��U�d���^~܈�������,���dA�>.R��s:`�a�(���!�zh��^V ])>~ô�8z�x5ٷ�&g�}�g[�(������M�:�E�(���|�3�YM��M"��eV�Fxz'k�Udm�������ٝ�=lOUm�:�p`g�t�D��x6��*��F.�-k] y�-_���JBvT�WcN��9��a�B?<���e�#�^KC1I| c�p�Ƕ]�������o�vې9��ROd��W���"��<#���EOJ�V|b9��ޘ�Gc- ��ҩ��M+�t�%��Or��%'����'�D57��z�[��(�B)$=����^���4U��~�D.c.gy=����Z�/u��Yp�(Ȗ�	�tmg��������Imǂ7x� � ���G�8�`�ۣk2�K\�FhF�ʙ�x�*����-[�����ZgJ�h�7�Nyƪqm?a���(~�}Ϛ���t'�Q˚t��[q��<<{s�/g2Ua,줅���|�|��I,�͛���&�f� ��:;��o|
��,���@�e��E~�IXM�G��{�&�ޝL�i�m䩃�0�7~��`���e�;�H"e\��}�Ӥ�N�_����g����+5���ʳ�]����J䍓x�!@��C���;�tFX��^�AV�d�2V f',o[����iD��C����m�I~��>�p�g�\�<�����Rm����k��
��g��$�OZ]
��~U�Kb�)�m��Z�e����n�גӠ�w#Bi|U�������!�����@���r � �L�M���h������N�������3��s�A�^�k=3a ���	�ۿ��)>��&�_����oy5�Ьۣ�ڻe�kKUA�1n[༤�<���>����	熮˳����J7H�0j����K7��lܽK%5�v��NFlW�5x��<]2PVф	Z��HP��Jsߒ<��|�pǻR&p���Y�@�}A�/�釙���x��*c�)�s���;; [*?���+��zs��/?�Jun{���1}=���1\�6����m��{
�b�U�x�:�7�C@����
fN�6��G�e��������W�hi{�)�%$��)�y]�`��|�#]3Fo�<s��b:T��J��V�)�k�˧e-�gK��[A�ߍ�1N>��W~��{TN����1�.�C;�Q�C:���c�F�#S�j�^���r��<:=�_ϯ*�k�~?�g��'�I
 mj=���O���m��F#b}ζ^�g�s�3n�9c�Tp�w@��G|�@B+����H�c+^6_�_H%H.��H�h�ݝ�h�V[��[z�},��Uy��8LNHڣ��}�#��X��r�P@���a�5[�3���E���ĭr�K6J�k�
�������fe9"��;w���X�&U��W_:y�����_bMR<4:���3I$�`OAꦛ������[7(׹��>�9ؼ��\9�*U�u�Ĺ�7H] =��L9�C�Dv)�-ڪF3��y�:���B���9���Oŝ�R9�ۣPU9ʭ�s�J���wf*����h�NP����ꥤX��O�$o�W��,�VccΚ� �hg@����|Lۤ����'��ǻ�ï���uۃ�&vM*��tU�:0��ɔ��T��j<o�R��w&9����nɻ��U=�E�H�d�m�s�r�	��L�=�h�hة������[�Q9�,�1�a� |�6&�f6����@݄�x� ����z��nN"�ߛ,��/�ˢ�������h��^�x�
$�L� ��#U ��&f ;�む��@5�I�9�6xus�W��� �ɀ4�
�\�����&A���7q�	Z�J�eOW
�@�<n4�'����-f�"s���x���ߒl/3��\ch��k}�>&|.q�#��FT��!�Io��խ�e<
Q�l�"�wj��Ҕu�� {�2V��y��A+{�B�n�9��|�;l�3Y�d<�2����g��Nw���3�#������Q"���"a���T���L�* _�����;bw�o;t��/,f�)%�v��)�g��� ���7꜄MpJ
e���0�\�!���)у�S��L�n���3V�����{����\��g0������RP����~��w�mfߝ�_��� �ٞ�Q�U�Ǆ��p��2�/�{g��ag�^rhA���ҟ@��pcR���@ws�`��~�W�p��9!�ǳ�i�z�x(3���������}J�\V`;��wƢ�l����OcL��� �;QJ)�'r��_0�=N��pNx�r�?^�Ú�pK�J l������dNT@`��_�ҽ-��˶�Q�I���!�'�kH\�3��^���wbq�uZ���9Q�;��9g��D�Ɨ�i�oI-��	�������>�p.��M��,��4�Td�������0��2�|ma/zKJ���c��[�m[#��@"�����1��HA��< �*�����s6=^Qo�*�^r��jEj�ϓy4�)��A�����s�a��[�ȷMxJL�t"��A4�|mb��R�
���i�Y�\���a��7���?�}�K�K3�����$l�5�"7��/m��J� d,��dǇ�{W�d�?!�����:mޟhP�JǇHn�Xc`���(�!�B�-v�X:,��:���u����l�o�
��Y#6`��\�暷~��^(4���Z~�Z�9�p��Hҩ�n���;W�My2����zv�N�]l�q�K!�|eu�e
:�����5:s2���D�oʎ���.��V��@˯
���a�Qi�м���P븭}����7>� oWu�n�����.��8�� ?�}OӴg���G�My�a���_ �]����}�1��J��*�� X&Enq�ղ���g�},�F�(��Bt���|bs*Z���|G�X�L��Qi��ƵX���^�QV��bq�qn=P�.��kK�5-��^��pMB�0T��9��S�zD�b��e�C��S�oT=�� ,ɂ����j��o��kٸ+?(��M��k-a���qW�.��N#i�b��q��]&���Z�$��r��๩m���`n�W�p��1/�>ȋ2g�� �����%H%�%q�sDQ	�܁Gxp������0X�A��b��KߞH$Dhy�-"V�oڼ�췛��݌��qC/[�Ip���
%Д�A�2���N�����.�K��#�M��XN�a�R�Lwh$���m��ʉX����Z�m��T��]���7�eW`��J�4��4��Դk7�:�.�Z����*��ƹ�v ������3�~G���L4s�z�ҸLo�B@ki.��a�ǜ�倞.���ө��ӯT�8V��*�ٚoR8I�O��>	��X������q�?���5v4l�*�?Cک�)��2rj����&�����#�a��N�F F|�*u�'����<�w�[�~��o2�(�ɢ5�:�qx��v�{G��͆X��7w��L׸8Y�Y�<�` �w)���O4:��pMe/��*z@Z�:��n�xN2u]���8m��Kf044�t]�)����P[��Y�?s�l�q�TgA��B�f^��� hY����m��o?�Ƥs-�����g��d[�/b�|�20���|�6�G�:i�(�ݢo`��1�P= �4X�[E�TE]�� �-�E�+-���]�Zi�⍻ˆ��ӕ�<.;*�Y�d_D��k����0�9��ڇ�WE�,ۮ�*�����
x�ȟ~�o{��re���<�ij�\�@���J57��	�Js�����Ɂi��&C9)C�^����|h�/�HF�r�G9{1�,y0{#��y!�t .�Y��	�=m��*�aܣ)RT_:*\V�iӊ�R}������ C4�-4���U�<B��F���L�OUL3�pl]���Տr�eݪc��y?��\�a k��n�kk��P���Z��!#CM��Y2��E&��h�Lw�u�=VY�C�������f�zR��Įv7�����uǊu���>�j�&��"H�M{w$.�߂n��M�KT�Kն��r�W�A򟅪�4�r;�Kg$yW@A (X^l��4ȺS���E�)��;ԓ�hJ��le
���$��9۫"!���y�#�ф��5n��b�Y٭�ᆩO��v��,y��������!���%V;����1F���0�!��]��+�:6��M���W��C�R�%ER���NY�	ؠ����Y��@��#nq���R��ґ�~x���	�N�x��%�	}��IEHB<	�r����]\�Ddضr������W6񑥿�o��
�+�l��H�j�. ������$P�̬-���!.C�~�
7R��U	t�j������hLb�H���x@2[Hwtx��|��S��k#$�S��	Ԇ�),p�]7�]��TZ�5�_q�����Aó�pG("g�+�_-C�*v�Ht]�Z�0���VŜ����<��J����{̗��I�k��F��>���'I�8�e��$�]��ԁ|��+��s��ģ8S� u3���F���?��%8�>�
��F�$�0�P~���I�+��+�;��R�QzK�$����1 �r�H�:>2ܛ�M��*�	�n���xW��䵽]4���ܣ��Z�(��aNAָ�7,-A�w|����!G]C��
1�<Y�)�����������3j��˘��8�X'��jخ��}��Zի�k������e&p�	�����MR���ZhB͂xӺ���N? E��](��L)�(���x!&=S�<E ,Wٓm1�%V�1��^�� c�2>$���~��n�Ɖ�v�	ĮK�� Xƶ/#�Hm˜�����[���?��{�y<˒����u�󔥾��m�mi�5��D#���S���2İ�^�ϳطP�=�ڸ���;,�DA�I���%�quD��v���)����j�D�$݃�������/��_f.���r�b$ф��Y��[ڪ2�=cWD�窃U$Fzd𐴑�� ���9<�(S&�bN�SsAUm�8P�,�G�m��Ǉ,�[w�� m"��ϡti��o��ɄD����97�_̛��qУ���)/�b K�.g���F���;����YR2���"�:���n�i��d?������Q�!�1kN���/���<�Dğ��CS�b+�\.{nUٱ�#�"�Ƽ�B��Z�@o�e�6S^$@�ܬ�=r 1���ąS]���kS��3�
��Bc�i�o�����z�Ѧ�C���k�J%'�T5����R��+֍@õ{�o�@��/����~޼�Ew���ƴ�j4�Y/�b�}G�l�Ⱦ�d)l1iS��g�}Q[���\�z�L��a�v��W߻���R�F�O�VXc��'4#�{����<⃅x�]��;�%_u�)dgN=tl�4S�[�8M�	�A�En�-�i�խ� k�Ҭׯ	��&?�H�����;5�w{,��Z��l 3�Pzmac��r��o�&�<�V��j?����%�{`ߞw�C$%�?������x��
5�n4����ZM�f b.�]�(9�LF��o�v(ƚ5�h��z�b��W옧�6�{��ؒJ����$F3��U#�9K��,�֐�h�����^s��O�k6��	Th��oCt��Ihձ�Լ�d֞1%！T�>��@����ٲg�Z���:�/�8�b��j~�ܾ�1�슚a���_�0/M)������y�|�
�ۚ�e\�{*%45d�S�G�;��v��.�A�����)���Y�Z�R\-�h��� (	��hu��l�F����:lЭi�b��˘!)+�@�u`��W���;����^�����i�:D�މ*�۸�\�E�����e�w�?�Ոs��.�@��H��JlD������Z�I��5���{��b*>X�\�
����Y/ �"��ɋ���I�cԺ��\�> 2mV���ĺ2"��ƀcO��yR��iZvc4�-��;�����Y��@�)������˩�#(���lH#uw�Ua�%��r7�L{p��ɺ�\jmd�qo�@��Y�E�wYS�����aT�ۊ��B�_廀�Y
�f�OqI�=�y ��������Ō�5=E����@ǻ�:��x�Z�7��CPm���b�L��]���"Q��'��A�Es0��#�p�������\@ϫS�D��f&���f��u�2x�c�~R�i�v�z.����ڃ-�}�{2�6�f'��C��b��^��df�5+W��3&1,]$���A~��4?q��u�q���J?݈��ʱ�~�b�`g�{w/���0���N͈��_�_O��":���� $���O˝�M�W4��Æ�A�v$�<�6x���*�]z������<��"��L��Mo��7��8,b���ܗ,)�(1���w��Th�S�x��[3�]��a[��5��M�)���`�h594 @Hߺ�JI޼��HBhPU����#�����m����_ �C��U���踖ak��I��QT�����5��~�_��o?b�C��=��$,�'2Δ���	���֙G���hyw����t�og�?0�1�O93�^?�	�6=��BY/�|>	���nD۽��rR�(�vk�=���k�(ѳ�H[]����<�
Xx���%��&�`�X����x��-Я��ۺ;�`+������+>-�\�6c1�T��7��k�@)�Pu���g�������ߑ�4 �~jy ������,�;��C�1��3?���� h�1��n�dsCܮܱ_�U��ǭF~0�G.��Yv* ,�z=д�l�>�����@t@>�Ƨ�fl\�	q��s8�X�3N.�Շ�z�`�9��g�H�����������+J5���������v��6���S��%�݃�xE���+<�9|���5d���w9�2�-�c��\��1���g#0�Dw��8���$uHz�{��J6 sFIJ ���ןB�$2F�B�����q+�2��nb�<�8u��7t.u	tg�24�{v�l0�	
G�l�Rt#���I{�$�ɁٰW�M����'蔷�*��3cT{7G���l����º��$l�9�~"g�_��rZ�g����M��܄�z6�=~ja�'��P<\���ڟ��������}(�"�҇��3e�ͮ��$�k,�j���7�/Z��m�i�ur#�q��`?\_����L|:RW#¦�k��H�%��m%ve��Cc.,Af�B���S��ɼT���g�f�����|�x�ĺ�ƫ-=��zCl����@�id@!l�l��Q<�������cL��*��{R?�ݿ,.:��p�Sљ�&P:�u�dj���<��/����#X.K��U��v�ǁ
Ws�*������ �/���nfD�-K�?��Z�y��'�'�nP��G�΢\�-�w��5�a��\<�ȶ�`h����"8�1�?�j�Ơ_��P���)wzi㸄{�2�p��c@U�w� �ſ������e��l7�ra��k$3P��iAn�M�x�?F׫�$��=S�?g?��</`��bam��6D�Db ��.���g�E��^q�D�3�f����l,'�=���"��T��O;MQaѦhܼ����g�PE��`�\��xcg�W���|'����
�5m�J����}2��MK����#2?�s9(����l�P��8��,�.��k����0����;v8�����|2��]۟��<+6�n0^��0��柔yo�%��Sݠ����#!ºo�g�0��4uI��~�|x�i�%�����]�Gh�z���XP&���ec|~�A[C�L^�N��݊hkf�y���y:����>x� ��*f
	�%Tk�뺘�mDC�68OH�}��r�HIj� �"�9kA0���s'�5������^��Q�8��#C4�ʺ����eɀ�6&W�qlqG�dq�)c��9'��]Ǉ�_�f�{4ȗެD�a�%�j)�o�=��F��i!�����A� �Ι�{п�|�&�]&k��)z?�4�w�u�DUS�  `I	GO2��8`��M&Vr����Ѹ��Z{l>����Y�j�����
���٢���� �9u�N�A�&��TV7��ߚ<�uڳ�tU"m!�Qŧ�p�U��މ�J�k�}U1a����bjz}3T��=_p�E�d���!O�
\p�~��m�g��T.T��V��"Z�n�:�H��I'�Ȟ�(?o�|��7&�qϒY�G=�Ϯ�\oD�fM�Y��4:���>oG�|CEu�&�K|�v�y��z�ܾ���a�#q���` ��V�}Vi*����Z?�Q`���z�t�Dgŉ��\:I���� .x�� ܫ+	>��t�M'�?���4����n:��9����D�kѷPഥ��ݛ��y%_cp7�|m�$g����߾�أ������"�g���EĊӫ[���������S����Yki�Bh�|&��l��Ne�Ʈ�R�]�4_�$���ZcU0	�b?�x���n
/�낷�r6�Nm��L����B�8������b��`��h�%�@��p�⋳�w��7�?��{$V@~�[,p��V�/�uopz1j��&�N��m�5鑊��L��������x�͹.�h(��H k��7��C��1��/r1G���N
���QB*ĭc�a	���9��]��Yd�l*�+r��L���%�?������"a�ꋝ�̾qkY)1��� ��%�?u��k6}[m���r�s<�Z������v����UXU`���M♀N�A��	�|7���YH��[N<Q�m!|��!��ɡ�F[S�ۊӣ���͡p���g33[�s	V=�A[>d����;��&م�,�VA�+�� ʒ�;}�2!��z�~��K��a!�N�.�����#����
�+��Z�MoA�S�K�}�F��:~1�'�X0+,�K���K� e�|N��ZV��(�����]ݥ��`t����J��ԯH�"+�,�0�l�p����+�3~�Q؝U�'𬦶X����Ж啫�	[�
�mh�]Pj	Q6��)8�)qCQA�6� ����6o�f�Zr>���!Ò��������a���ᇝ������� )@��
���8wۉ�勢H� ̖��di=��|Xt��࿛�`��r��o�uG$g�ϯ�C�qq(}�_k]7Ǝ�@��5����U��m��Ӥ��]�śѸ����[e�xK8ӌ�.�`qtFb���xU�q�~FSok:v�,Y�
?%����c?98H��L���`����ҫ���П�G��{w��;-�qB;X�4Q��z{�,?�2w������3{�r��7\��ɴ1���y��9@�i�Z?�T��n�g
��k���qO�fã�Q����
�tp��ޘuo*�CvIm���V�6Н��e��Έ3��:a�Qm��*дs>�9{�Jx���.�g��¤?�{���.{e�+X6��8W����{��eC��]������Gw��l�8�h^5�ać�U?X��6%�_$����#��Φ�����{��؞�1xzG�X�n�%N�B��Q�2h���a������kL�29�"�[��.�n)���ӆdQ��:���ك����Tt弛��g� �!�>���ec��R�Ӊ'S9�����h��O�Y��ƃ��������A�c�P<� �������dui�����5k:?��h�k+�Mvuni�� ��#+Z=�gk%��޺�[�*і�X6|m��{$Nn���ۘ��l�e=�U���Ÿ��+��T0/g�:�al��ؿ<-�=���ֹL�����'��F��)�� �WH�k�N�E����F�h3�0��Oϖ�F3�ǈ,p��$����|�.3*��Ȁ��D�tp�'����s;�h�1@�c��"O�� �Zo[j�u�}���w�&w�:�B�H�����Ў�4�\9��̼���Y0��ٰ(�����1�����:���7�Xڄ�ޡ�����Xޡ�E���+Ibg�)����(8�1�������<��}?s���S�xalӬm顛�7N���Z0�}�$(�����@A�����"�����
>��K�^?Y�
����J�۠�(Yc�󕡽�`�'���#,<��wN�x�v���8OiG��}���Э5��3��r��\D�띩"��!�wE��pt�J��x%R>\R��&-m�k÷UD��
��5��H6�>� ����MM�i�Q�D��-�/@�j��l����Z=�q6��&S�-�U�T���G����'���6��k�t`� 䥻���/5f��#>�љ�d������t�bJL�\r����d9Fb�A5^$�0��E�"R��c.�S�K7_`Ns��5�9*�6,\[��5\m��C�%���ڎ�pŒv�ח�2J�K�lhC��}篈���z��L��kj�r<������Pw��O!F;K
�$P?�@�ԃo�<�m��O���+�l���i�G���5ZԄ򝤒��Y�:�c�� �d��sߠ�\wUD�";(�u��k3��@���rR
�
�c��c'�Zr�*�3�!��<��TF����L6Ӎ6m^04��J��&�	t��g�c_���B*�ua���qɞ�eD�%����bR�Sf�/^/��?7h3��/���CQ��~4�>%Uڳ(+{O_�CL�Y�5P��}�
4�c�o�9��ΰ��l5�~��4r��C�H]%*��N�m�C���\�+��'1��J������.<�Fd�II <P��������_�~���p<EI�[�~&���N���nσ�(K�</�����/G�JxՁ##3v���w���:<����h�b�+�Z�������7�(�z-eCl��gzF�y���ח�}�&��8VĘ���߆&.�������.�9#� ֏�ao^���9n`��2��� c^�zP����D�ў,���@:���ƌ&���5�H,�4������S�	�+n�bx��}�0K'���Ց���Uf�.�m��f���(�g� >��2�W~��i�o��ߎJu������<�X�>k�v�I�c#��gs����Hbk�_���p��c)*����^�}�IMY�[�)�M����\�gaz��*yF>� ��X����m�|	&Q�hm �
XCD��PE�}ʬT����0%H��:	 ׶��b�Vx�
�V+�x<ba=S�T9���qwt-7��=��ܨ����̗���@����?_K�W�7���zĔD6jS!b���� ��2S��o�5�_v�f�>	;#HΊr��9{�! E `�2�&܂DOzT�d��4��F1�vˠ!���wcJ�?4���ŋռ��_|)�r���[??l�L�7��	�ڋ�36�K)��/��sq ]1�Uv�o��o�g�e��۷�q�Gp���< O�~��Ek0g��� (LEQrNsu %�y-�g�u�|I���wYS����>k�����[/	�f�T��;&�\l���E�*h���,��_�)�W`d�
,P�[��N"rx�ht�x�a�tr|����ա�ۢ��2�:�LC�#\V?]�O}I�/)��o��~��#���������=�ED,�C�����6,2\�zs~���w܊��-�+{��$!��G�����c�4����Pu\j���s~,�Ou�Hfn�(�	�u8��`�b�<G��>	[�(}��>>�F�d��ϕ�~lfMmA�d�E�ĆUHC�'o����lO���2\Y�~��R���Q9D�t�7��>l8���-�a���	љ���Ov�[zO,aO�˿�u��p�|Rs('�x���$G����<���r,� b(��67ӖE<]������MO�Z�뮧��}�"��o�,�G���a��4*s4���6)Q�M\��2+��פּ!���c�=�?�����A�]2p&���	�l��F6�����[T��w��#D]�������`��27���ioT��(��������ݏ��<���a��&�ʊo��ܩǾ�8LA�����ԛw(n:���z��A^�}�fz^�����(����7�$)E��A1J�8j|k�x�u�B-�F�z#�-�W�(!�f�@K>Q͕	�j_�_-U)��K�J�6^��w��βr�m���̓����j`������cCjW�$??��g[O�Z��������p�?��Cl?�o�io�V��ms|<��2�]�kuy��|�B�PT��������k���g�GME'���j �������L;%=��1o���ƕe�O��f�.���w46�rK�.1��g36I\x-rv�7#�X�@��(6ȱ�!sO@� K�z�W�Żw�܉��5�sj�_�ep�������,��V!�s���@��2#G��(����"�f������D�P |��uX��_�jS���vѱ���	���S����_�hr�y���2Y���|�qDB%�7l����#�S�c�1��;����/ 8�ɳk� I�)M����N���3�W^|%����]�����"A�GcM5��:��4@�����6�-;Tr�q��@^&���+inelK���L�]0h�JO�}��)Zw�/��l6@[U�e��0T�H��^2<��ŀ�
(I��b�����C(����(��l��P���Q�LaE�9�D�?I��W�d\��8�?�Q�w�������=����g�zO���͟K���5;]�o-�Ԇ�5lh�:N.�u9Ϩ��֔<���]4n_�� ��A�>D�VyɎ1b��	_��f�}��Gb��V�N~S�3�zLb�w�S	�Y*�]��
{xs��vH�k���]<U�
m��h�%�1�Tkm�5�o�:N�p�7z������2(��܉:p�.c�������@�$X8���p��@ۙ�j$D���>�<��v_l.R�]����(Egl���y9�>���䔝�B�m��O�ڇ~(���R#:Yc��*�������D��t��N�#׻v���b �,r��92MFp,! � �`�F`"P�y��v.�XڂՅ���;��n�>8-��n�80j:��E�C����T�&fO��N��_8���?S���?�$1���LE�zX���B@��Y�\�Q��QG-�;��Ԩ��SP)��^��Ţ����Z���V������kNr=I�c���,���;�֑1'خK0l��@L��n����/LJ�D(M*���]E��H��J�RsnH�@l�]kBB�<5In{�����gɪ���x4�/�@~��`U7�q���Yv�׾B6�G���	��t#�3����[�Y��R�s{�V;r�L ����,	r#Zw��ξ��9�#���0xG�sƵ��R��2\��p�D�4��6��*���s,V���u�3dײjPdO��MDI�;�us���
\����ig�0?@��Wz�1W�E�*�6�2	�*���Y��L�ס�D�
�3�J��~;N�e��l��
��{���:r��(;k��x$����mBP��v����Z[VT�@/; ���j��+])�z��Ƒ��?Ea�^�y9׎�����D �Q���M`���۔��K��V�FK�{�U԰�n����"t���Qe�6�2��v�����@O(�Sq?�.�?�5a}��K��:��i�(7z���(���A�����N(N:_����M�����#����p��v|��|=J?�!f*k�Й�]�yIY$:�.'�3�0^A.��}1��Mx4T�5N�(?=sH ����.ɐr���&�E��;VEA�9H���!������D�/�_}���'�J�:z������`Q�� ���;p�~;�C���-B����L	2)�vBa6�ۼ�S �L��.����$�9�f"Ug���O,N�Y)= ��9�J���8C�F��VrLfl��P{l��	e/��J�V�� B�}�f� `%�����6�ʚ�陵<<:�	#r|�/̡5'��V�R�ȵH�A+��_c�LT�>��zP�dz���)x5_�?�n����''�{���;��jc��j�t�;4��g��>���'M[3�z�A���EZ�Q��on$�K��p�]D�4yQ�b�8�r z}Acli3L�L�羽�H��RJ+x�~�,�w�Q#���JZG��XÇ��Y�N�VZ]��xE��Z_\cg��G�#�����j,�0� zr*��;�z h�uF\��dL��Lt��<�0��c�a 5�K��Ho��o]Q�؈{=6���帷����eD|¤��i���W`,��wMo�sx��S'��1BK	�F幛��ߚ�h/��ܵ�ǈ����.��ܹ��;��o�1�����p=�)��r��Y9J��wam0�������r&i[�+>�?���[o:���w��<Zr��M�*C@G��w��y�9�=�������q6�*&�dv��
y�kW܎��T����q�.�C��c����U�d�B0��۪�����B����;[o�M��=b6V�k��
i������U���^� ��� Fs�W%��_�\. �A�w��N�q�>vΟٷ �~8(��SMe�(X^ǳ6�c��o�7�|�iQ�W߻z`�k��>�ks�ހxǏͅ���e���d'�Ca5L��э7�����t��M7R��5j���'Rna�Ƽ�Q�^�RVfS8��R��
��<�pkb�SV��cN�:g&etH�?s��^���=�V�k��@<@���F�8�Å��7sw���.��o�*b��4fUt�mJ�Ʉ��J��x���YU�O�P���h3ZVEq]x�����/��9� 7*K�FLJ++�Ɠ���+�QB��'��v��"w^IJ
�V�']C8��(�Z߲fa�.��(N�,��>!9#��$���^4��T�e�<^[T��EU�cۀӯN�c���	8Ê�&���@� �Dw.���gV�wUTW�B]��+ G/0@-����_�!mg@�i�7�4�P���"z��U��(��	���t!��|��}�G!������d�\|���6�t�m} �u��2P��Nh���ePޕ|���ld�fpa�b�"��(���[!�BRڟD,3�#ꍍ�I��sԯb8)��z;�3���Ǜ�7�WL���!��u*ro(�ܠ5�&�^��A�-�G���}����!Z��[_�&�*�A\��[v6����w���S�w`B���^�\���M��	�ct�a�~���T�'�"��}��o���#(�B3��fMv��}�Q!����p)~/Tբi���k��C��.�����ƌ/��x}��r���;��z�mB4tR�&U�(�-Eލo��������{�-j}m�$��LK2�}�D�s��)�{s���u���^wIޅ#���nWe��LƻӈH�\ֽ����'u���'|tmZrPg{&����R�L��V
L�x�V�'W��-��u�j��O?j�ߠ&�j|���h1H5'K��He%�bȠjTsta�5v�u�g���_
0��R����B-�0&�[�4�~��y,��q���W��T,>�{��Y^�Q/Ã��ȉ��C�*��ez"�m��ͻ��O�SfP��S�Es�u.�N��KN���dv3+�ty�/�f*0W�ԊV�{��d[M�}����^}��k1��;/68ɃC����V&?+���ŷ����v��㈛,^�"��ń�~� �����.P]�h�8QE����ձ���qz(�.i98y潴���`���ע�C��/@XS�mUm���҂K5�(�+�E�6�Pb ��79X� ��5e��kr#���F�����n�]��yjVM��X�P��j;���ʛ��8�*�I��W��y�]�#�`���4b��N�F� C<�Ʃ�|����	��9}�&ށ[��f��-�q$A����^�/�Յ��ix�`a�)�-*:���Y�W|6����@DA:��%�E�z<��T�v6� �b}z8U,�ڠ���@g����9�Z.&0����ڬ�g/~�<r��3��˯���=k3D%�0��9*ىd���<ֲR;�^҅�$#��-�{�\�*�VV�ߢ���$�~�jy}���dp�������;2+o� =�],K�@�KY^7@���	�W�Jb�v��T�3�����6W2������6��"u������^��U��#�K�^��"����k��?�%&b��������'D�V����D��_z<F�o�)0/����2}b��݃b��d��6���?�s��X�c�*H)��1S�B~�
��GX�t-v7�/�W�<���!X \�%��(9pW?�^��Y~���~k۝x�PQW}T�"�?��;y�5,t`�tYSq���F�Z�p�	�W�a*83�r�������*���-1�<���y��Q��6�GDP�bT��DI}pN��!��S��ݢXu�j�O�8$uQ)����F�������:�2����sb�W�kK�1T��KLz9Z�#�W��ӝ1{�q�pY3.�S�c*����,�����M�?`���	����I�S�QH�uoa�B����V9	A</�m���\��Hr�3����=�q���(�fvUMI�#*�Q�"��V;td}ʋ���:B}N�u��D?�A�Jvc�v�ԨG�X.���oK�m|�^9(���²�cF]�!LxZt�1M��\$�0d�YN���ݣ^D�D��:!wy��c��C��5V�64�&����a���t�6����z��OR8�h����E~oV�m:4������'7�:��x@'�rZ�s�:�h�9c��	���ƫ>@!�r�X4��M���.[�R�8N7�av�����W�dKf����Ǆ�<S��D�pFFU*z+�gT�@G{$&Ê�fq�lYl����<g�����9�.@���S�'�E�`Po�"l.��"ҡ�=� +$����v������^��O�4���Xԑoα.M���e����)3��j{�o�:|���NǕ�7G�v@UBpB��<^H�Fq8��Z�
���,��1�׮�?=��ܑNa��}T�;����<zx�]�[�'��A� ��p���0��Ԃ�s�c��Z5���u���f��Ϳ��2d�6XwI�����m@���D?:��*�~ �@٬�v�Zn�$�_0��=J3/Ʈ��{�8
���d�������P����g*nᛁ#����4�&�Px�|����K�� ��4�����ӷ�	�G\���{��?U���v�o-9˶�ڧ����t�"(+�_��>�\������r�̘7�S�Պ��'!?>��Hד��Q���S�O~G���o}/&�>QS�@�XS)vV�E��f�����QX���Ȋ�r�j#Ώ_�S�kazd#��O��J%\T��-E��th�|���g�ș��D��Z-�7޻�ҷX=�B����6�ك���䦣Y��4�	��r�M��|jN�����q x��'x���,��g�~c�>h�
�)�T��ڵߘ�����.E!�͘es�<���z߶BM�Ȗƒ��(]�K�M���p�Cr��[������w}��\��I�Yt���/7K��v��S��q��m2����WQ�3�wA��>�g|�5��5���&̓q�+�	�NN�޺q*v��͉�q��\�i/$A�����z?a�=]]������4�g������˧QkU$�V?�pڦ?w��މ8�x�>5�D�O=	��z	hQ)v��~=��gݙ*�bׅؓ�m<���g���3"=���y�˱�pei�hl��)���	o�9捍]:�M19�)z��93����O�m�]��hei���7�D��]�y���~�q�^Ͷ��`7���Ҥ�>�������	\��+-ʕ�Y���;W��PwMe�9���
C��M�q�P��~�(��#�/��9s�Ȱ]-�fIt��k���Ṑ#�� 1K!��!}�#t��cW��|��9��rbHK;ˣW�
ٰހ����y�na�K���<=�l"e��*�j3����A��b�"�;��OK�LU�R��I��ٹ@���к�PH���>�U軄4?�5�H����̞HbM;�f���Y��$8"�v��\yĬ���c�Ю�/��[HT��	���嫿 � :M���iHr{�Qy��D(��y�W!"/\����0:D��Y�PN}~ߌ�K�l�<#
��p7��i:��)�(�t��y�K�hN����gQfIc��V㟼L1R���P.�����,$ѻB����~#��Jat��<�!�� �J�a0��FAk���B�@7��u��]uov����S�Z5C����5m��ʧ�l�^�P�?�_���Kc�Q�;,!|���US���	��2�p~���{�`��ݯQ@���E!t����< w_�n8��_�"&9�wcsu¯�+{E���#ZcU���Ǎv�
�S�/��P��$G12���uh*@�J4� ���V����CWY�`�`��l9���ూ]Ȣv_����t����V5�jC�V��j��6	A,C8�x�3�eO���΃��mGq�.!���|b�6uU�9���|~Ljw��|�=C���V�K�	Jg���� i
�f������0�0c������M�y4��cra��zw�A��ʀ�\��}��5U���M����*+�#�}��xy�ƨY�Yn�{���lb�k���!��QC+
r�#��]�5��j�^�)z���8#_�o\�%~��D��`zL&�l�[I�%����N�.�".a^��|�S�ӕ�إ�����1d����~��Y��1��1�^ǆ��y��dPF&j:���T%2k�-Gn�^���.��W�g/CZ�M梑Bg�l8�e�6c������x���6�����|������aՎ����q|OaS��<���K�H"�,�rm�kd�Ǽ^���8 v`9��9�p�HЊI�
�Ck�Ӄ��G�kڨlUٚ����N5�Wo6=�Z��,=�^2t/y��:���7�3ͭ3��9~�rY�}Z�)���F��0��ݷW`�6��/�K�J�c�ԯ�Z���O��܂Κ��!�01O�߆�q�����so�gIpH���2�Sf��:���r>N��ĵ����� Ւd��|����\��2��&���ԃ�xCt��T۷Śb��b���e�����'��"�и���� �o�g�}n/�<A9$ {�V�.$���)����ذ�	��" ���I���Ⱥ#�4��;Yb���
�SD����L!v��ߢ����
�Vs=u��i�8��u� �R�1a] �81�p�]-.���[
�g<�&$B����C[CM�,I}�lƊ&���O@)���"I:t��u�w���=�`�!E���z;��)�~��L�23�q�ͫ�8w�!�ĝ�je�xFւ���>�.�兎��\���食}$*>�a�?7�Ob�}���?��9��� |�5�Tf����������/|8�@� � :C���g�I �B?䇵xC���o	d��ar����g'|��]3�Y���!A�8�DI�JH`��_�\�Ѵ�T+�N���G�i�Ζ�X�b$�?��<��U8{��hm����{�&(<G����y�����<H2�� ��]��G��&w�2����`��̡�Uշxޭ�D�8��'�:(m4�!l�q����N(�eBxX�Y4�� 3�o�{I��1T�𓊥&�=aЪ�R�Il�&ZP[��xe�Xg;��Y��a��3�$l|O�Pc��(� *�!K�%&OO2��#V���f\�#a��x��=!�Gw�h6gv�k�͗�mf��)jUu��h��4���V�J��լI��9�N�W��ROQ����H'h�"�ہ���i�g�R���M����@5����B*W-Lnp�ʭ�@��i��+[�g�+I�]r:��r9"<����fb�Lp���j��I���z�a�Ԉ:���j��ܦ��p)ҍ*)DU����fJ}^�@��X7��]���R��VOј�Z��{��3Y3'�]1w:먿d�;�1��^ł����ۦ,e�6��)JB�2y�����O�4�Y�RJO�Ś)@���~P �	�h�SnL���Q�`h�\H'��iJ�N;vS������[��}&7* iq=@|�6�@���q^��G��T%����T��*ԣ�
��
�,j@:�����l}7��?-��惂$M��m��&8�w͝E@�j� x��*اk���b`z��q�ՆnZ�F����b���Ţ��wX�F������GD�j�����"nIH>ӰO��'4�%P����hT�����96��y�¶o|�A�[�J��?D�H<%'�ND�䇻��� ��=���4���^��>��5�u�8�B�Z�;�=j�0�]JhoAW_$�9���g \���W�ʖ\��h��F�"�s��}�Sgѫ}md���t��0�.��]e�0�oZr4����
I�euك�b�k)RL��uX���M����u�,gJ0��h�fcp)��	�:���K��+~�ѫ�ie�Ýɷ��D�hry��Æ�Gu�ٹ��ާ��XXQ-$H�Cڏ�E�<~e�ϱ(��)�פZ�EjN?��r%I`[�KHw�ޭt{e��H�!e���V/�DA�M�N���%:)�NE�`a��cR1�-��c������	u���A̅����N�e�3"�
��v��T�{Ƭ���_���%jc�PZ����n�Q���̃�)n��Zqk(��j�a�I�1��_�H�jG�87��e�dGz�G?hmv�4�A��`<���ۍ�?|l�4B��`@<1�1�z:�z�v�wV���v�����ez�Q�B+�R)��&�Cn��]y�uc�0a$SlĄJ����MR���q���.��1?Y��)���DW�����$AC�V��s�P�v����H0��0��O�޺J<�/��j0�7+=�������.ټE��)p�&B��!t~c��y��f���p�d�o9�{�A�x��]`�^���#��^}��yA��.�|ڽsf�l7����y2���Q~%'*�w��~JD��{�[����v�]���0�@���o�n���B9������e���2:͑ �yGS����ͻs���l{����<�g��Jt
�Þ�V`��6�#�>���֖X;����a�S�~!o�o��% B�@�А��C���D�X��ov�kSx]I*�2/� ��ko��p�M�_�l@����Є��zI�.xy,ww04���X؂#��^Ea3�h��ҏ��r���b�x��y���{[�{<4=R�n�/�yQqہⲣ<ހ[N�%��	ȑ)�xQU�_��oæ�  ��"�Z�{4�I��,�n1�N����B4(��bX!$�$�#�{*WTFB�ͤ�]���T�K�8+�^YW$q���@�sk�QS�Ҳr�q�&����-��FZ߯S����mo�[,��D�P>Kk� �~�j��v���N4�3���x����n\��gTǷ����z1n�p��8bG�>T��2X��Y�C8�i���j���Qg~�(	!��k?L*נ�!N�ep�jK�Ic���F�H�6������q�D�шr�������`�X���QL���� z���OXۺ�!���zҹ�[�b�k�l����6,W
?���? �Gi���U�H�G�&`e��.��>I�e5ihj.�VK���
YO�З��m�|ׂ�I��W�(,�]�2lQ����H{����e֓��t�~4xԫ\��-38%��vj�)1�i�+$E�9���1��M���=�n�x�h���:�5���'�n�"�����6�^w�AsI�ű7P�Č�ֹ�7ٛ;���ٛ�9,5���D����S�683L�hr�8��@߫@�X�n��17�, v���u9�j�K�5h[��]c��D?��St����W��՚�ߎ/�����`O���� �����eU��~R�
�Z�*��59�2��.C}o��)����a\&l�fG�Wm{��Q�D2�_>�µ�
�[AIܗ@�>Ť��WI�hٗ�J$��/�q< �A	��PY�k'�Wm$�GJ���X�O���)���f�ȉ�����:=�δY�ԀG-G�G�X	�[M��T� �w���S�V8]Fi"�R>ݶ��.XxEH%)����v��5m���Әv���[a�X��f5 �%�ؼF�i��v�~��#Κ�P�k·�3�0Ğ���R
�ıO��/D�o�<��,�P�Y$@��U�N]�ZD��Rbx�-I@���]����Q�ǹ[��R����42�+E9��8S<>)=@�
�P��ݤ�j<G�����V�=^2p��uR���/�<D�f��nY֯0�@S���ᄾkoA�����@����nA����@K3{��v����� �}�꾵w8y �Bg���b�)�JP���>@+JG��+
�Iæ#���|�;w�&D�`voF,����M�U�����k�|�*{����P��`e�Q�fd��;>k$�1����)���&IN�/X��ԫoh&�����<t���a�+B>cC;��|2���6��C±2��yO�&�U�'_FQ��u�٪��J�}4�Ge����Ot�_Ƒ�G�A^��q͆���b{�38D���T��Ao�\���L�P��l�g��W����4Сq�Uy�81���m�||�ы!�Z��������Ȧ�p�'*)�_OCEA���3�k3蔨7��O������v��N�6BuS�q*a=�q��G�����^685]�z}O����o�ѳ��6�Clx�W��~���%��j�\�[��<
$ɏ��X��=(���[ �5Jԏ���io$;�$���yF�����aY
�1��R�V,4:�����;�-AO�H�����:��+[�h�]V�\�U�T���t�{��^į�e�O� ��TVx-W���tT�	'V������V�n�GPT�&��W�_�J�֤\
9[�v��۳�]��m/�1�c��������+�5wuo�k�y�҃W ����M����_Cv~�B��/3�0��a`
'�T��Hw�&3����J�%�L� �i�W9f����m����Os2�]�J*��SDc-�5�p"G�@���:�5�c���TW���8f۹7�=Q��-d�,�z�� .��'8�q6��e�?��4~ (p�d�W�����<�)Zɵ���e�G��|_)jmj�>��wv[��|S�\�}�
�f �K�ʲ�ڇ������^T&{��)&S#pd�c��!�+I ];���p�5�S%n��|�L(���|w!{��e����r�Eꃅ��5���K	yx����Sv��O[W������{b��X=ۺVo��ÀFݢ�s.X�;pqSS�b���gܒ�C*�u��ҝV�< B��@�'��D|wc��p�����Di�b�#C=�z��Ml��x�/�d�V�!:����T[�et�K~~k����q+ 3!^��Mٚ&����.bz{�$7��_*2�
��s��Ӯ2	;2Z�/Y,k���*2%��0��v	32�"(2C~'`K:���s����~p����D+�Ma���lx~�P��tn�[s���Ԛ�,&����|*�θ���.Hk��z������ln�e�M߼`�LʶǞ!�_lR����rԲ�xL�x����/���`e��\f�㨮�8[�Z_ȫq����5���d#Q9�Pi]�-|�M�/[A��!l����~6HC�{���M���pm�9��/m�Y2��x�r�=�T���	�%��4y�:�*M�u��>�;�G~5u��!6�<+W ~>$�Re�[���r��&���(���/�q�c��y�\`Vn~f�sdWf�F&��^�2�ޕ�
�����o�.ؑ3/;���U��Փw�z�� 엩;�H�d�g����!� �&>0%qF��8�dS��5}��Q�D�:��B�+���9�g��w��[��L(� ��7��ׅLJ��J��$�<�~�:쏱|4��]�9/�`5� K�kLl�-������<�&m�~���`��B됲��d����,S��v��͉d;˳�轋�p�PU$��-�!�,��VP�v\XI'����:�.�%"N�at�A��e��4�٭��IA�'����PÈB�o�m���+PX'&�+0Xb<p-ف�79T�Kz���_ൟ�Ov�`2��6̨A5Z�E��Ͳ�g� �d܁��E��sXe���nт�d�@���95�ը~�8�Gx����
�9�~9P�gbP4�����d�󁋇�h\]��wzуm�f�DSk�A���T�f�{^�$�]Zw���c;)��9u!^6�-�����(����r���B���`Ex
��j&�i�󻟛ƿ��[v��W�UiU[��u|���/�
�)^C뫋!tbP�n����#�땫�qu��0	�vA4BJ"��_Qn��+Q��W�D'?��w����>p��(��/�RXF�@���|���rwpp��S�3ؙ�T6�%�e�YY�D�U���P�Aw�N�_u����/Ko�Q> ����F��x�Y�ċZ !l�j&�|�`�����P��ұƈ�����������O�3[(L�ń�g>��G�+�@��]Vg\��r�by9�_j8w��������F�������(�4���=�C�y�Ձ2��1���=m�D�$px�71�}�K���>*͸|O���������=%>���#��ӆ�c�o��v����_�+�kT�G�L�L.J>�;B�c�*���KK-����M�۞j�,�ͥ9�U�p��n����M+�����R�,�/����:`[�bZ�L�!�qY`��~��Q}��b3/��70��L�G
��ch~�/��0ȃ�jB*"�ג$.��5M�z�NX���X��E&ڞ	W�.-n|*�	E&q%��(ٺσ]{)&���@��Wj=E�B�*F��f��NPiP��xz���7��ӥZR�F����-�gep��%h��$K����[����@+�T0��F��J��{YJ�Jn�{j�K��)�/��	F��t�c�w�uB>����X	�����Tp���O%�Ҹ�!�f�l"	]�F���R�ȼ�l���ܑ��(�?�\o�� �[I���3��n��\�Pp�_^� ~yI ��$���)�/��ͅ\���5v`F�4��8��QwҦ̴r9
T60��ɘk�	�l��a;@I5��W�"y��Icw��E?��f���<��,G������y��/r3Pd�3}��%D��!��V�-�u�3��Z
P���PV=��u�j���P���e����G+��'H8]�N��wk�-T� (����`��`���^��9���yAi����V���I����4�>c�Z,B�#��T���K�t㧕�5�¼�Z��@a����J��2<�y��`��!	Y�J�+��j�.�Q��ɪ�٧�g���M[�@�t]�q�aeS�i��"�˔Ӑ����dp�E5VI,0��1���fLӥM�:V�w$҃S�U��8�|˅G�ro����EV�0j#���w
X�{����A%1���|�ŭ�z�s�BU"Nl

t�A1�MB�O�K�@o�W� �K�C�Ɲ��$�9�f&7��r��Rmװ�����I[��3�V#���.�ߝ�	9l�����.�k�Y`�&,F�{ k��&�2��]]�ؓ�g%ߨ$�'-%i�t!�������pC�������B�1|ԙ%K��=������(Y �&����`��v��B 2��e/8�7�uF捚Ϊ��E����pNaeҡ���"Ŋ4c������R��?��cm�F'����*�r#�5,,w:+HPg�E�<@���ݸ�ģ�]��P)V>1H�e��R�ز�<�3�d��ֶ�
v�`��ۨf��PYAz���1�wʉ@�d:&AlN���5A�('�,8L5AY��[~�vn<I8����כ�>o9�K���"�57ڧ|��vsoT�.����G5QPk�	;��úF�v0�N�!��>�����W,�r����B���"�vȃ�X��APYvʎ���uD�-N+d��قG��]����Y�VO[z�8�@5�;�A<���-B�5T] 
�"D�:��WR� G_�����z7v�M ��&���x��4b$����A{�>bu󒕠Ԗ�S��e���_��M��Dᘀ;U4����e]������La�~�G��2�Pߎ�m�o��1��:�Q��p��X*Z�Bx/���`�������	�6�/��^�O�1�}�.�[lK0���:L�n�ջ|a�k�Z'Xh�"�;�R��Z���MP8|�x2U��-+�h����C�C�s-�6��Qh�$z���3:*P��K]���B��x������ۦ����G}2��k�@�8$
�}�c*%'��\SF����:��~Sl��|��UE�T�%�S2�oQD���Y1	l *9��`�Ɗ1����HK�����r����FX���!AqC�#f�w~��0��zFό�D�f7��v�:��|h8�֛��;:1�B>�Z�դ�w�	3�nmN�����N�-��e�J�ڮ�]w*����D�A��!Z�m���p
5����o�}��ނ�������>ъ�̡	����lfm�qR��i�"'of��x�%���hI���8�g��V"�<&� �+AG	 Kg��iX!a���R?(g�$3�	*2���ᙹ��۽��FT�2?�ی���ڏT�8E���5g�9��27�QQ o!Dˍ���PƮi�evC4�=�f�qZ#H���@E����I��W3Hpo�����bl[�`�K����N��u��+������o�)��{a� �$�$���T��|)�Y &[|:��a��Ήӣl~Gk5�.t��mWa^���>{��t�uolE\��"���9�==�6)^˩����xp��S���p��A�QuXrX���VB�%֯ϗ������Y�+}b�wc��IȖr? ?lce�T��8!^7�^�%l��p�x�S�$@�_��i�x=����S6��o��=�}�d���'|�uH�*�ز(8���mܮ�:�������	C� �גVpLף���݁'�ɇl��}��*�$�0�T��8=}hz	����]HJP'i�Ѥ�ɪ���k�t=��U�KS` �G��I�ձ���P(��詢4¼s�$_3ΓL��+��ڰҎ{V��ŚA�J5"�X�I�'�b��	�]���K_�������'r�+���2�Jz��:
r�?���F����(D�N���d�ם4L����#�B��ݏ6�e���U�EFB=����E�K(tզ��}����/��x_�DR��:�I��j'���;�|��7�m��)�k�KM6��m��)ځxL�1�/?H"Q�X!:8�t`��&�'�PuU\�ao����vr��V�hT��ާ�u�����`��]�@�Xǂ3�OJ(��N�U.�h��Rc�#c�R!6ܘd����e���R���r�al+��$3��Ƅ���n����p��d�:;�xi̛����"���n;ʯ�j�!	�a� �ٱ��0��ũ��q�ɺ����@�`��A�6��Ȱ��Z\Al�v��������V�` 	yk�0���Eٹ8�*�������$�		���5��.8����pnR������LI������u]�P|�_R��q����B� �4���:����.dv�QH�ɐa꾈�3� �3of!���.0��1�׼���8.�s�EB�pئV����PS:c��
�fPc�fqx����� ��S�2��8'���y3����)H����*�o���D�3,����@����iMP���g�{��[h� Vi��?�7�e��6]^�B��i�YL��A��Zȭ��h[n ���$eG�~x�*Hxd"B�����f�HJV'!���xr���'~'X}8J�^�0�W~_bD'��kgĞ��j}|.!*��%R�Џ��3�͟��о�K�׾���]�s+��|�1���٧s�Y�f�V��H���G*��P�)��4�m�z}���c���d�����~��6g�Ո?��f�a+p�ԏa���}���r��lvm�<�Vk�֫y�B�&_	!�s�@��L���"�y��߃۲]� 䤮��m���jM�0������=7����qV��?�y�R�=DO�#�=��4`z�e-�7{�w̞�:�6(�T��oem��"zK[�V�@i���_c�	�p,u�V����F���<��eFv�I����ڋ�Ko�v�Yt�MP&���~�q�еO�޷�����|v1x���@�O͙���|���Qp����)��|���(��.j�js�[ȃ�ik�D�|TF�o�xz��;��b�4��vۈ�P�bѺ测�li��������#0�E�8�=e�S�Z��M�w)�m9��X���	�Uٙ4Ut��LW?�
���a��0nG	����1�(��#�ߓTu[�1��&G!������S��ƭ�Կ�dB��sѮ�(�e���"�c�*�b���!��]*t�iq��W�5��'�zy��#� 2�!��w.��Ƀ�;�k)]_������j�F x�We��P�1~���'�Ң�����^"�2����Pr���h2l��g=N�c�H!�"��q�z{4���TWP*����7kgss�=�-�
O�ȥ��F�Jsb���KP��P:�5�Lu,��z�x����uIV=܍��8F��i���R8������X��rM�1o�㦓9��I�rLX�ޛ����ɵ�`]g�<�{pe�7�}IP�)š�T��QƀX����-A�;e��'U䡈z'>��nv�J�@�Έ�^hM��
+�[�A�V�%O-.� �Ѧ�e=}�-�ʅ��_���԰u�J�q����IV|�gE$HP�V�=��MHɗ��X�F3��f��{��+e��a�m:��8#όXD� �G ��P�_5���-����Ȩ��d2���
;*đp|ha0� e牉��T�7'�L�"�5I K��9���yM��h���g����[w@c�\��9��g5���g#�ء�哩3���hX`�I�f9i_@; ����g������,Ǔ�;�͑��t��D�uH����{����Fg*�N�G�5�sT���n�u􏹁8���.�E�Vw�LH#�Q�8F����)i�77�~vx`q��[�s��=S��q�4&N�0�`�Ouq�mC?X:�)vMd������ݽ��/l�zWGT�/���-��=����oI�!D�U=ۦ^.��u�h����)4�B=֬��g �����?iځ�����㚁{����1
�A*&��LNM\iC�m��}φ��+p�����S��������S%��d:��Բ���1���U�Ç�F1Đ���1�\�;����lAI$�w���\umPj�UG����f*�n�k.ȡL]h�����$ÓOp�݌/��
L6�}��l"����Nذ�c���iݓ�� rӍ+��h����㚞!�����M>�f=A#�`D��x�rz��%
C���/�k�RG\��@ج���)ԫݍ�t���םɽ���}�ʪ�m�R}�'��K$;y|	�=����TQ����ZB���+4�nW�G�,�^_��R0��8�m���*�䨅l;o��Hy|�	~ۺI�!�s����h��9Ee�Ԟ���!H� ��he!{�[p\_�Z�k�j~ns�@0��n��
�*f|y�r�`�)𝷈w���*0�.u`Q�}�mDL8OV�e�0l�ՐC��R�\3�吘�߫N[��F�&�S��+O#I�V��<:�w|0��m~7u��D���m����:���]2��2a��aH�)p(Čۂ)���s�JW�&�K�g%����i턅ɛŇOF�\1���m>�~7��?c\A[-R���3�]}�l��B�ܝ�%d�] ����u�0!(^���ɋް£&���6��s����G�!p7�$�@N�%v�L�0� �o3�(Ơ�<,�^77����q���x�+E!�)6^䌛֕T:��h�<|.	��ڮ 
S�>	�8j�a�/��r31������6�Sw�s��T��NM~o9�P.:�1X>�B	A�T����2)WS��9��~n���,�J�-�/��<@F`R�|�G|a\?	��c�)E�]��v��=@
˹ɯ�Q���'�)G����PHt�E�eM5��ʶē���$&�a��wٙ����J*�$󀮟l���Ȩ��|�pR7j�v����i��|���{��fD�l���e[A
bf�3"��E���Vd3]���� ��c��i� �8���,ip�l�Kd�
m���x���R����?����M�b@_O���L_���Yӧ�nw�<U#�E4b�ɿ�F��3gq�5�MH<���٫�٫��vjE0�D ��,f�u�J��ڷ�&/�J�%Y�AǙ��k��{؎y-P0�e`a��'�R��m��U[&A�ȧ}�ɣҎ���эl$�'I
���ܓ�A+tEM�r �o����U\|dU��1˧Nq��yS�P_"92�~iۛ���Xs(
�J����K�����[kj�!���o��fUŨ� ��' ���3. ��Xu(t�_����+��!jB*/,��xj����3)�����a�PQ�=y��`JU���Z�ce��Q1L</%Њ�P�;�ߪ]�}���<R�=C�ˇ��u��W�
��e����j	o�/G�./��{�{_���� S��k�1�x2����Ư���8��q靍�9A�ZA,�Τ�h!�N)
����QX���t>/ ����}@��
�7J�����Ҭ��V�Â�:s!�m�O�ۂ���4)%@q�9�v.,
���_�����[�-U�a��H�
}�
G��/��]�;���
���5]]i]W�$���ek�ǆ�p��A����q�)V9	��v�Y�4���H�߉�Cx��*`�-�h�2�%�j��,��k��X�Vh1�o:�(ֽ�\�\`R_C��ʹ��������b+O_��%�(�F�s���͉�:4q{���f�GD�K2��w����0�U�w�����B��z��q���x	�K%!I,j��x��#y��p�}}���N,y��_R8E-�_b\�HR/3̈�� W�ll.���+��m���X3�9
DW��k��Z��_�����?�H������]d��R�ڎ��(�:�|��!�D�b!���Q�(Y�^�}p�1V�歏*k��)W��_��$�Ig�����]R��sj��U�f��A�HTs0���L����z��Ncȩ���q=Em;��Yb0�V?��S�X�{�n�d�\Ҫ��AN!�MP���Pl����`~��p�d�<;ZX/1����4fh��(g񢅷�x��d��Ѻ�h�f<�Ӽ"
�y6\����O3N<Wt)���|�/w�xkĞ��l�[�wv��n�<�`�B�����LG�h�-��-�E�`�#pG;�	��,��#G�+?Dd���I|w2#�s�Z趝�����t��Ih��<auE�fX��fx�~��e����\������/���پ�zՏ@�̠h��8:9�"�?d��X���	��������?Oj��D����&�s�gZNqǊ���!S���$�x8t�GVc ��;�W�N���J��YX�C���>[�Jɬ� >����d�/4�Z��1R΄IHb�=�ƐA��� ���X|���$�����;Y
�\M����1e���{?~���2p��X/�Ǡ
<V�	;]��J(*Ą��yp�i��}UU�*'"��������Kc�u�Rx�ht��@Ӗ<��O���mk��`��:!Kq�^�CIsy�p��#yE��15WA Au>��jsq}d�-E����}P�$��Gj�䨇ܸ$�-ۥ�<"�hG�#b[�-[��DݤK���d� Kڷ��݌2�3f �hy"^%:�.n�{���>ˮ|��q��l����J(�j���6ɹ.��JEˇ<Qz.��0����]/DHr%0��9�_��@�����ד ���+�f?C�w���a�Oa ��¤��2m�cD��.�`�����`]lX����T^dR��DuKN��,G�	�F�����I�9L��A>��8����uU����j.w�\!�(]���~���L��"aĒ�8�B��[���W$jjcWV���`����e��6�XQ�2�*�Z��I���8U�D�O���:��O�6���F2�_����G1���y�gK����s����O��JW';��-���3@�IdPe��������3�.����������F��VZ��0��˄��;p@��,��u����'�u,�~�,���㽥\0��֓�t��A&>*>�S�o�/p��@o�dw�E�w;pq���5;my�13X��k����oW��HP�}�5�e8z�0�s���trI�۱\��@�6Gb����?~M`�܄(�UɄZ'R�'�I�u灝·��S�0q�Ps!����A#��b��9�U�n��t'�r���\�Rq��90���Ƅ��ҫ��5��T��%N�N��+���k��s�!P\�O0���cV�r�*�-l����==��9�W�B�,��XQ�2/Se�:�楊��w�J��V�[���������z�;�����;��j�fOf|ڒ�[���Y�C�YU��#.��I�ny�O1T�ј���8�^Xx��L��b��*����J��=h���4=m�p�b6�?�uo��f���p�W������.�::��՛�b����pӻ�����=�м٣]�3�i�?�o(��ɼE��n@��9<s ���	�
�<$���Xׁ��P��Qf)<}o��d������1���'��UqF�@�g���2��G�B"b��Mؙ��(���c�sw��]L�V.o.��\X�ʰ�����qV"	w�GG��.�7��Q�a�bwS�jA�q�K�~kM�܍�DZ����~�{����">('�6\6|;*m���Qi���J������l� ��'`�05�d�t`�J�B��'�@�e�����'Uo�D Rħ�X("W����*�ً9�K� )|s��l�ޙ-����8��e�X���
���>�d}�5�܃�����S��p@��DJuD*�O��Ϋ5�� �Na���f���8��勪=^����ъ��X�i��2�mt��1��ѽ��|9;�iE������PJ���6���b�d;-F�놘���$��҇Fo���+���>b`��ee
H �<����p���2�Cy�!9]���sD����빼����Ŭed)U�Q���ʩ �bP��8T�W�s��K�<ә���1�m�G?Ȅ�`��f��a��c���si�y���,+��'�H�)���/��s�n��έ�(*a�⸕����I><�~����į�%�4�j,��'��
�1%���Pw�ђSI���rs���iW/�t~��B�{��>EU���GK-ך/�M���IP�Ԯ����pFi[�i����s�I���O�&e���}�qzW��]q�T���ϛ
�I{ݎ�
���v�Ӈ�)���T�#.7З��/A:ތ�E���)���.l,_���r�K����H�1�	u�:=r=�'��.5��[ ��:�R�z �?h����ί��M�A�FB� �<���ތ_��woٻu�����4��Eh͓-W`{5\5 `����q��:��������-e����K�����؍i���[�e��t@�`�F͝n�"��Y��W���{����-z�����G�I;b@���u3�>Br�g�+n ���5�h�E�x����ȍ�D��;���?%/�68NTO��Okc�w>�l5AM*�8���>W8����7�@gg��Ƌ0��r$7h�����
��2w����<��`4�#!U�XxL⥷��;���pV���1��9���>�P���M�)p)s��uN7�0��6�B�:g�]U5�!kLIT��P�7��oy�-!i��(�/�Lm�i8�__��-�hU��?O��!7y��^����j��c����^ts��H�s��$H��&hġXիe�(���f�v_�#P7���`[²�O�ި��,l����cY��Xk��oU��Q�4L@�{B��r�|ܱ���l���Ď�mǙ��u�ڰ+^�-��fD�����_���`c��ӝ6�D�Q��j)y#v�l��'�bzD���3:�d�<�-<�r��*��<��Rk�Av�>0���f�#P��}�t�I��N'��1(&#7;#�����&����A!�T9ѯX�H�e@��8Iuo��uxje��4�ܒ9U�NS��.Y�t�q�}�#�B?��+�Mک���cC����(Z#���I�Y��u�I�8����U5�i������'΀�q�����GI��pw���g̈́s�����:�\�<�e�N�z6��5��U��AWX��^(�G��{g�[8�\����/��T X���G�f��>4�8+��ѳNq�9)�v��80ʞ�0�4*��Q�r�5S����Or���#C�>O�C����̢�I�� ����݈B�(Be�0�UĬ�hD6nE��g|��M�$lL�EL�ʖ�؏�%�{�3�>.X���E��  i��]w�Ԯ�Lp@AP��=fW�# �����M��^��mJ��ۻ�_��Ȼ�:��������"̳���;�ި;q�D��N��:9)	k(Y�ap$���MU��~��(m��r��#ᙲ:�6��/�

��ш�2P�'��s�0�*�KJkE������B\�X��.�B�s�R]&E������R�ʄ�H)�b���=����?�P<*ӝp)%����+g�O����
N�j�S�"���I��UJ��a��!�a� D&YJcA��\���Fuc$d��W��x�f���x�����9õ��!~mqP�A��pee�'%�^��NwthNѦ%�#hG�KX��{3�`@��_?X��+Ú�0�@�5ƍB�a@�RWץd�Z8��<;���WB�x����>�鍌WV0�
��ǒ�OS�c�b&|�R�����=')�O�{�1�;KZ1N�w&�.x�[�>���L�0���S������Q��/	�"�1�]+Ao3�y����B����a��ׄK�()J+��`O���J%�� �X.o�?��Y;��T�Ŵ��_bY��Oh���#�@E�сc�'
�tC1�"�����a=�z� �j���=xi:}H]9������
�Jg�Z�랑��c/�r��p��$9�ޯ�O�r�e�F��N��Ot�5����=�L�_�F��+��a��B���%a2�����4���Q}�o$�^���OX�+G��#�\{/A�c��r�_=���$�
��It��I`�J�a�mU�B��GW0�'��!���X�+����Q|�%���`��:}���>9Oat���Z �Vp?��:�$*_b����*mI���!�`��h��G�Z-�&�����}��X0O���|Q�M��]�\���BV:d�w�"0�"?��[g�_)���\����9�- 4��fN�Gjϋ	H������M��c��*Ĥ�6A�
B]��D�3x�d�0�����+#�M}��׆�?�t���EH�0��<x��N�{��Lq���A��0�~�htj��(V�����D�$��%��D�JV��^WzЬ��p���H��iw��K{.`��L�y)�Ӆ2ںhҺ�=PGr�nY�j������{�VE�Gd�=6���xJW5<�n�����uR�0AG~&���f��gv�S�s �'�e\B�Hv[M������g���5�X֘�;`�3I�0���t ���E����ū�1Ĺ��%K���j�C41=K���8I�ri~Q)�"+uM��P�O���iJU;Я�����pE�@|���{��
���)-��s#b��Ϳ~>YqU���2�M�wj�7&�3ϝS�,͒�#S��ұ��l っm���z��J����Z��s�?L޹V�����@����~d����������e��H|�w�e�KlŒt��e��,X���+��]�`�����Ο��b\��x��Q�$�4W��9���y\��(�J!("'�u�;J��k5��!�)g�*��y�{��Q��C� �zW�*�8����@6�h�[��`��R��X��-��a�4�u� ^P?���Ý�`� U��(�?�WGu J�LbZ3�4��뮮�ZZY���e)�V,8ȝt
�����'��d�.�����p��na��n1�f���t�n~�+̰�C���_�{bF	��ӗ�9!A}���D��#�$I69�Lf+�@ׂ�#�̂����>�O��8��@<��1&��������g���v�+9+j���u��>6���'�ڌ_�Y4��l��X��U*���z�9���Hj�,��|}ф���@��_�k��&�,�2�Z@j^X�j�2�`��dԇ�O�F�e SoP&k�V�`�H.���Z O�v�v$����2'�'���ဂ��<��ٺ�mϲ��s�����5سu�~n�yC�%8DeZ�v�z7y�I&`|k��)��9����ǖ�̱�F���#��n����٦\�k�1�t�62�[��s_�V�@�#�
�P��W�tvY�A'!�s�-=�#�K�'�G�&^�K��u�̎��_��;�`�k��4�<�Vw��;�Tm>Lۃ?��SE�u�>�0^#���:�%��|t�I�bž9.�8�<(�j��z>ήZ�b�[P.I�M
��� ��C�S�*��4u��&��vI�R�B�!\�ɕ�4�O�z�@F@B��a�AeKV�`��0HK�풙7���d��\W���Kl=��N��i5�qS��'�K�9�-
4|S�9X�d�S��[��3����@ۚ�� j�P���MWJ74h�}ζ���I����@�*&[2�.2q£�L�0t�ٲ��2����u�T^��>2U���v^޳�����[C�������	ϔr�� ���G�!�P=L,2�C�ga0��q�O�^� !+U��^�}�S��1zt�� �$�a��C�3���������L�&-"��o��lv:��p�W�X|��Pqoj�<p8����A�mI��J�77�s�,�uK�����"��ɍm)c֖�,]J�q�����g�������0МDJ��=X�aF�h��O����a	���Agq�R�12�
�'B$�֦]2Wg*hU"�-$tZGˆ���Z����ѷ��f#V�g5;�`t�`���ͻ%9��,%]���s߃�����p)��g��Y���Pr��	G)R-��\ �%T�KJ:ǁ��2��]�t4X�mxK�ꜥ"�����{�d�Ǹ$�Ɏwҋ�����
�Ɩ^�|��>�E�2RJ{7����UA;A�Vj*ns�6�)^��i����܆�Nƹ���n[f�+Ƥ��x��h�Ȁ�yqܗrѰ� � P7�s��.U�ؗ����֋�NBQxv$���R����}����'�O��gQ�O�/M�p��(� �D�3�FBFuۊ� ɏ��xEd��ߡ��ܛ�R,o"p+��r�����k`�Pc��]�^��V&�ر����d��֞Y�$����%7�8��wU��n�	Wy=V��`�((ǌ����}.���[���B�otH���7�;&�ON��(��3ue�NK�\$). ��_������奻��4j����5�����|��R�FO��_Y2�xZ�m�b�@���?y�,���Nq��v��k&�.�ͱ�Ѝ{O��@��fE��8�2$O��.�j�/�czV�Jz�� Ծi{k&ih�l]TBb�jZ��/�Hs�B�;0��QnE=_�}vE�-��޼�p������l4N��d�^��?e|hͮ1�)�[9��9��̠(ծX���*�o ]��2���0;�z��;٥΁��*<����.ۅ ��63��&�<�Ij��6Z���NT�M�@�Cb����{���f��+GG$�L��އ*��<aq���c�{Lvj?������ �z�:Itox�%�����.�ߛ���&�m�"es��T��!�+D�����
`��-���޻HG��}����!dT���?Vo�i��F����Iwr���2g��;'�@Bx"q���v}[��mu8�}�eN{�= lqc毈�r����6UFj�C�7�qeZ�'�\�ݘ��`�:j�� �@�}����%��0�v{89
^A�C��W�ʦ�C��{�\��l^rW���jT �PVͧ�];	W�1$a�>FD��
��z������H @C�������D�w�*� �5f��ƚ� �3��1
<EW�ɯ2�*R���*-����d�����c�b�q	;��T�c%K|!�T�S�7IK�1I�����1�&(`.2GC�!뢖B���"?����?���C"�NV˙����Z#���4��:�9 Ԡ-0��ΐZj�BQX\��@���?�WC�|�S%2��� ��y��G���@-&�1�}�0}{�΋��l���-� Y��
�&�lPo龐Ui��ҟ� -(u�~�b��WI�T���y7=)���A7��}��s��@�����>��!h�V\�kͷE�=���g��9��( ����*�m��w�>��ޏ�o� K�������Y��N���1�`��$���*!JUޚ�/lu���c�9�)�䇥��q�&�]+�=�*�$TRڬ�H׎��/r�*;{�H�cM�c�<gH���eT����8J�9�[eD�%��9c�<����$����~ǥ�̷�@�{�A��F�Ưb�j"p�xM�<�ͩ�!����o�aH����:��}�ɛYRlc#�}������a�_\o���D�#t��}V�����N�>jI�X�F��Bb���ƿ}��j~��G�&�Y���AZ�V�@��,_���'�oNo��4cZ�IH}y���C�/oqH�t1?8�d��$���ny'4���@�F��q����`����65~�kz��%8�_�����^(�y�F���]A�qI�m ��!��M���jc�p��0�3C��M�.X� 8�q��~���Nt�`!��h�2��� \k/��.��P��ݙ���xI�%��i'����+�R�����7-ԟ낯�?�P{R (��ͬJ\��`ۚP :h��e������m�9�/L�H��&�oI�Z��>-|Ҁe�ءE{��Ė_�_�B���ސYJC+n^�<{]D��? �� s�{������Q��v':����QZ��uM��4�w��ɣ-i8m��r��K�y� %�R�M��8b�AIh��O����\�;r�n�����"Nx���o�}����?=�yd<d��O���ă�w�C��+������'���E��ɣh�9�8���=4�9wp1��W���"��J��_=V@oU�v��(7o�_^wo��^Fhaܖb����rT��r��RP�3���`@��ʹQ��ih�#:6����X)2��n~f�b��U�]�R���EH���1w\�2|)���-b��Ӛ0c�KP��*�/Ve)��g+��v~���}8b��EW8�&k�9��u?3����s�ny�vQ�;�Ri��)��U��g=Nk';��mlJ����FrZ-�sCJѮY���Y /�������9�D��X��>
�?h��E��X�A�S����E_Is��t�$I�C	\�_i�(y��\��6���=0\)E�%auKք�G�Q�&�l��u���4P�4j�o6%D#$<NlX��*��2]*�����4��$�>Sf:������D�A���l��$hE`漿㰹�(����p�n���"�9G�Kb!�j���riVT�%а�E�4�$��S�(��,�ç�ߓ�v��~k!}��A7<#���"��t%S��iW7&-��VkM��<�w櫖��.���u��Z0&�$+C�u�fC�&ɤr�h�3?�Ž�0�tC��`^��R�kp��v�F�?��m\+\jc���eXVDdO#�~	?���_�`�y�|<�TͻNnw�Wݲ���lW��)j��C��L�՛ 1� =S��-�[�1��h�h���_�I(:�[�h�(l�Q,��ֵ��)m�I>i�I8�Vu�����?�,�S��7 S��*�{!�;����t/� {M��k5%�Gȏ�9<�	��^���#Ni�^���0y�1�BxaɡdJ���ХfU8W�[Ip��i��;��2��D�e�EhO!�>�e����bߚ��G��<(6i��f(���v�4wƍ=^(X������ʑDլ9�4��� �HEr�Uc�h�Nf��~�MM��H�/QpA�N7���9>~�]Y�{���R�;�s�4Fa@:'G���9:�:��G���)=w����Q�[��w˟�Sg> ��m�z?�C�5~����d9Ϸۇ�a@�1��&�����γ��+y���b�-A���XJ�,8�;i���vJ���*�$Qm,�ʦH\�1M��l��1׵��#[�ߴ�����L�DW.���ЉV��7��ݚ#��Fa�*
����	�(�O�֜R~���PG����i��F�o�A,��zzŅ��}�#��[���3����\_�+<�~�*������Z�y��cЅ�9p�~���a��T"H]c)���^m��<�˨�5�	'��
��n[�;z�� ���!ٴ���輜C�.i���N�/%t{ŋ�����9*�P	�6��9���?D��y�@�,�D�����<�h.;��*T\M�W�O9�Z�8	,�+�Dz[�+7!��,��4��yT�#�0,�0��Eq`�_�Z��|:�C&�?�$�ř���F��_��\8�E*���������Q30�G��Et`�@��$1٬~/g��֯�� U���`0�W�?T�{y�}�ә�]]y~��EB��y�e����Z�E7�r�%s��k�Xb�����M="lr8!����1���dwS�r�g��y�Xs����^��;������1&��<��ˉ9m�{�A���=�(G���e�ۃJV�:U��/|^I�1G���'�faz�ɢ�=91,��wJ��QOD�6�@{h!ϖiCtj�E瞵'y�ah5/��Ku�w�"���F��<Hk���r0, �vf�x�o=�Ӕ�"�6�×����b�l���!nx��g�Y���Fǧ�Z��K�B��$�%�`�u[�=�Ao/e���t�$�t%��m�䅩ͩ�!���=��=�]�;4�o�Cd�^X�퀎^����;vm�Ւ��E�D1��� ���`�C�.�jy`��h�3����3�+�<1+#ۘ�xM�a���^��V�Y9Gנ�c|�pP��n�_���'���>�5�l�؆��L�5� �ׅ�YL��Xb�~Y[�{���v@�M�dэM7Z�M�γYq�p@H�-Ѐ!=��H썄)������qV&�~�e#�MʂmZ���'�5$1'����%���p>?��R<�3D�T=����&�X6���$�����9a�A@ 0�,��l0��sO+�[W��3����t����_@���/�5ʼ�?<J ���j���JBG}4�����?8T8(V�����8"ˋ���MTC�������uP����8L/�|��E�I�UӥH���~f։~r;C��8o4��E�/�)���.l�q<��?�j����w�dNQ���T-�({�
%eݲ�~!�F���{IwL���t�OT�i�(J�Ƌ�j��@�����&��Q�G�%���!����s�|��'��8��6ƿ�� cG����p<>��&c+�4a����(N�.߲M�FFK#ID@��iB=�� ;%��.�)H�^:��Q���hZW,�0�ڠ�r�%R��	��S@ur-3 6܏|��7o+:k���� k��T��6-�s�W@��T1��$��Fh��C��Rل�.��z]�
���q�G
��4�ݟ*&+鷎�"��\�϶� A�e1�q�<>`��J�`�LJg�pӹT��Xw�uK�1�MZ�+k�^#�i��]�6�q����1%w����W��P�a�ڒ^@[�G2�+��|\E����lLB!W4������M�N�\�f���{&�\�nd�GOР��:�"٘� ��(�챃���we;��5�~���Y��c���h�7�v��}/���^�M2Ǉ�u,�r>���5a�1�3��Uy�Ih���P���W��EB�ˁ����0<��4�ù�b(\��f�bmC}�=_�H�[�U����2���bd ]��55S�l=Lw6�EL;ju�n~��i�$������a{�bo����n>�)��/��_s��2̴���M�5�k!����-#�㏔u;?%�Vz,�S�S�sI��@�I��=�u�`���j/�בA��<$���$NC�a�gj����z��s��V�^��m��V�+��v������h�8Z��`���������S�}k~�`x��§�?ߧ
�5b�ǧ5��2>��F���gğ	5Ě|nq�s��gcvñ<ހܪ���:h>���&="w 쒰$]'>��2����J�&A��w��4J�⒘�w��5���e芁�m���]��޺G&<X\ f�9�,�}]*'Uݶ;����������싸���}߶�t�7w�6�Z�ϲsl��ͥJ:E;$�U�zu'W�Fcg�����jv�3�����5
��?{�Bm=�:�x�-V�'Q�cݱWoH�����h��n�l��I��e�̴;�<�LjS�%�݉�T���:����>mo�"=�[�.d���-lQn�ժB������fr}"��]<����f;&	�E�SJ���4��dt�f�eZ�'p�Nkx����H	�A�֝3��׫���oH�I�3���YU��L�"�`2�4]�z�BN>��A;PpQ��%��H����|.��i�Z5������H@a�Kt�@+y�̦)�2i�H|�e��u/Kj�C�>���,�~��3.������x������^u��X�6Jќt�;��a����g���s`p�w�P�j6�#P8�uh�У!��Zc�fճ�����F�?�SZj��E�B4?5���2U˛b����z�+��mE��j0�v�Ax7���~-�#����H�5�������N6���w���`��G���c[��tt6v�ۀ��^ȲWW,g~���]O�<�~�#KJ����]�E�:�K�������x	��\��y����R�3��q�S���=̓l���U�0,��1'0�k�A2���=�r�bfp��y�m7@�0�H��^��z)���{?LD�9��t��5kƵu|�8����j��5�ͼ�ǚ�a�5��w��@�d��dA�(�Ӯ�v�v-u�`
ň����[X�pW+]�fYY0�k!��Aų�G���D��:�Z�Pș;n[?QN��;����#kG�4o�( ��kY��aF(�w��F�Q2ӯ+�'c�Wo��C	��{W9J������p�0n��Z����8�Eˢ���h7�f ܩu�y9aP�F �"Ӌ \G���Ż����TY]�r��f��d��P�|u����P���>ˮ�1�[gP�y�sj��T�l��B���sr��C��m��E��J�|8��zj����"�b��<Pg�	�t�������\��I�,77\�����������M�0*,d�T��\����,��,^B��闘lyv{���
Θζ�*l�v)�)h���D(A"����ɬn���ү"�0<�[S%H0�-?�����/�B����D��A�D:�3��%���IG$�q�h���ȳ����Hj�^v�y\r���6���߲Z��k����f��t�\�T�Yl���)%x�n�C�ü��Y�s��2����%qkBbbڔ`C���;�b%��O��B�������;@nU����q�&��x�U��-��I��֘1w�i����W#��
��"�=
m�G�����`k��c���V���:�?o`��R�1K�G����Í3���O�!^j��;/�f�ԓ��v~��}����{���	��k�id��`3ʡ^CkJgO���g�;5�훗�@�s��R'�I6|�Zz)�=���ǒP��XM������sy��!�����Y��S��Rb@o����`�8=p$!
��S-�v9��;3��'8p:������A%��ڒT&mg;��_�1+o�b��b�}�}녗��|��x����Lэm.�Q���r��X!���j�~"�W�ޢ
	e��v)�q���*l�_�j�W����2�:$��b*�h]>��	mY ��g��PO^N$9�&;-iAj��<�xW���9��ʑ�'�͘8t��c
�Wġ���HTU0�×u0����O��v?��s6���g����X�\�&"y��*'�pU��Q�p��]A@��\�~,�2`A:��Q��B~�e��w@J��,�*ɖ�-�{3w�Ջ^�V.��ͥ��t��+�b��V�2ls��O���BW�DD?�F���\/�dIL-���pA!u�VH��WXn����\:�}%�L�;���}"�@��v.2<��4Ϧ�V�G9�]����n�Kew�QPN��$-�ۘh٘����ʼ�����	�` ��8u^��
��KG;Ux��S�j"չ�k����W�E���a��X~�)�� jk� �wX�sL"fc�pF�ΐ�� 0r����8KFt:߄p��߉�,�~p���6��$A<_6:}����j�] 2��>��,4�����X��c����r�^rs���� ��n�-h�蕫�)+j�����m��|�!{)`�H�
J�z2�����gWzۖ�*8�EO����"�����H�3�0ml����9��퀺���[��Ίc�|��a��vZ3թ$@��g���J:~akl��M�k96��g	{����t���c���Lw=r�8\H��K��s+���k ��� VK4����.�쁷�r��}5k "PR�8�D����&8Iy�J�|u�t���{T$�Y�WW����q�zs���\���2SH���`��0����]��������3���u����g���p��������z�<1���'xZ�o��N���4��o��D̛�V����wTƙwRV�i0��ڃu�_�O�]t'�2�2�_���D&i�'Cm��BELĺI/�py��L�W2���ǉ��BVy�������̃-t���f�#-n���P&�!՗�4���q/�\�k���O�N<�P��lF'�u١ȥ]����Хވe�O*>)-�M_���� 8�A�xg��#�n�2����;��yqBF\8�s��p��;;'l���_���(1���愃	]<���K���[W�s\E�z�[�}Ъ73F�$.������n�Itc?��i~M�`�s�л��� u����:.��2SI�$U�sR}fe7�p����.��y�Q�t���G��/���˶"��~)�+�P	q��
��+>�Z>�;֩��m���U�i�N��N���~���#�F�,�K���	����%(M��$�:jvݑ���1��-���3%�}����Rpk���7㱵�hp����6���ƎM��/ml�D��fnK�P��]���NjP����v�ek�2*3��s%��W`�L�r�"�+U7�9��!	Զ�"���!abfW�H�m�����j1�r�����?���8�?*B��z�sF�����B�Ȣ�i�fb�����VV��s�X����џ �5^ڸ��x�{�иB�(jh���%���)�x[\�:�ߴ��gm;�0��Q�:|5ݥ}��2^�M���7i�!��~�k^9����CR�S�(���u��bM�1>�Ζ���G���%�+�wP,|J��p4֟�x�0�Ml��=zq��d-�9K,���>�7�6Vꮿ�C��}�ʰ�oV�O%2W�(D
��ָ˷_����s�ၗX����1�FFn�|�z����,WO�"�(�&�l����W��h"w��=�Q�m��g��w�U�>u��������[�7Ϙ?�����Ȉ���ɗ����w�8���)�����p{,>6֍@��=�\��JAb��I�#��� s�gay���t:R�MeH��Ã����Rog�y��V��Аr!��mՓ�dU �{;ȑb�q|ɺk�;��}-v���,|C�
~�^j)P��X%�l{�~
�#aw������G�Q�!+}ö�@ѩ·�Gl��FC������:]�Js�� �5���[;��VU�C�8}���-�A����}d��Ǣ����|����9S�>�n�����xE1A<�k���P��M��D"V�嶽���k�����7��q!xʊ
y�ud����pj.5[h��7��b@�^7�lѵ�A��I��J~�����U��3\�j���}�팊�>����]���B紊``�y<�n.CY��e_$�1����#�O�N��8}t����T��`UplصwzN:�~��n��`7�� hd���+L�A��# J��S�U��_��1���J�Usz�^�B����y�LU%@0�蝴s��Ea< ��D���.��>M��Q��$-�\(=/(���dіq��x�1��k�~�le��QIiu�h&�"�<�1I��-��Î��^[�=Y�b��~����ʼ(3 y��ɤ�qv��=�'�(4��Կ7��8l���u�~����
�YJ ����n ��+Wz+�XV^�s-a! ��t!���˲�(ug�![ ��޴�Y��-��0W@����m7DMni�~3O����@=��\#,��/�G���"�P�:_�U-_+=���ήt�<���W����J��v5��!�߶m��R�K���a��0��]9���M������}���6�EbJI䀿=s*3_^�d����1Q˭�&��Whi%�fØ΀�FhE�T�RM�(Φ�U�r?����4y�JW����}��JE�ւ>OuAE�o�5��~�JZ; B�Sݸ��on|���Y�ŕ//f�C�F�O�5[�fG�s'��(�J�8ǡ�Y7�_{ܩnq�^B䘹�Z���zΖ�E8&ѧŪ�K��GO��eRc�� 6D�
W����o���-��A���?s)B� ��j3�6Hh�\�uQ����YY�n��Tkύ8~��D_�Y��,i'8%Y^dN.;W�[��r�� �t���,���B(2aD!���K���//�&s�@�[͎5��������5KD�鵫F���a"P�,����ˉ:�Nk��r#��\��?p?P�Br'�K-���s��p�H�2���V0�+N	���r�$��-7����
�]�д�^�>Ҏz�o�����~9y�ɶ��T��D
��>0��Ι;��3OÀD��|����3˖y�|��e�[�vy�ͻ1���-�;7.��F��#��c���Lp��<nfX�H�:<$�J�3o�W���D5��#j�^%�䬺 �,�1�\� ָ!�R��>��?����Rn�'9���L�(:�
N�"y�:�Y����[u 4���0�4����b,�A /:����2i�Ų �Q��h��חJ-!XfU4�O��=\7�	o ����q>}���#S����O6ܲa�䣊�ap%�ʊZ��8GwϽ�Y���z�0�/�l��0	��?cmY�DE��Zw太^��o��#k�1��w��JC>�L��"�kޝ1�e�_���~`�t�$��$��{+h2��~�[K%W�����*ѝU}�075��y���/��nD"�����!KG�u1l�:�X:�ߺ�8#�}�郈p6@�?0��R���{�;��k�+�,y��Q>8��~x�[�4 BXX{�o�M���c�0�=:��w�n��G�u9e���4�u@�y�c�QMS�z��l]�8��ӌ��q^{ыῠLi,�V�(5-]we{U&7r8B��CL�7����4"�;�o��K ���3I�5�#�]�Z!l8�1*�[+�Q�5�&�+�**�[�z%xv8�ؕ�?��}J:�;MLBWj�����h;������0��q����FHJ�\��i��~�^@��Rg�(oTDj!�n�	�<>����N�u�U�T�V��M(��ן(-�Jɧ��n�T�*T���B�(�$BUɘ��gk��R��!������h��5����Y���8+۪��ߪ�C5(c,B���؀���R����o���1��,.Ǎs �����:q��~#<9U�b���I#׼{H<xO�daD\��'G�et �I���Vi�Yi���/s��ݕ�J+�����\��a�R%%Mh��.�G,���
��
<o'�0���v�5����=�e�X�0}#�!�%�����H�v(�R�"��]��=[����=��}��<�v���ݚ����uq|M��SI(,�_�8f��q�9<����K���B�{�t\S�d�:i��BȞ*:w��xF��g,g��G4��zf��5��o��m9�_	���p�z}����WCz~[#��C훊=���[c���k#��؄����D��#VD?����D�}��r� �9v3&=��w�\Sz[u_�uÂs��"���G�_�+Pv>`���4��	W�7���yg'F.�L��h�Ddᨡu��,!������p%e��@�q�����!�b�닄�ewFY��9�x4ބ�ƥ��At�h�|C]�G���K��[.VN�ٝ�Vg3k'��q8����9Ýpց�%Ň��Y�fIE�MQ��n���%�n�T�ʉ&i<�D�U�Q�Q��k���i([L^a�Z�� ���:?�{�X0����ct��k��=`��ǀ�[��B]�|ɝ@�sq���[%�]�NZ̥��04%�������
bf#�T"��c�XР��ZY�/�j��.OM�u��ɨ����&^290{�r�Q�KQ�7w��[�,^�z�����C���S6@>�,,=�#�Ԙ��L�4P�����e ��t�k�����_`oG8��%���	�� �1�d'/;n��n�=�ä�s�e5nIg�`|گ]x�淹lʻ���u�p�j�	J�T��6Ԍ5���2ͳ��g���k�`0��X�|4���f����w7/�Y:�R�o@}�"�]t����j����>Ӣ,���C�2P��
!`��̼[�~Q�DTRd��-0���0Ӱ�AӜb���Y�D*�@&��r)��.q�=�m��( �%H�H��z���Rx�F�D��P�>Gq��D�H�-#q�V*�xj�JSC'�����a��n�og���.Ԍ�i���v�Mi�*zQ�D�8�T���^Q�͙�,�	2g����:Vπύq������:y�l�v9L�[�B:i~�,�_v��X}�uU�d-+ַP���yiec=(��p-�0!(\��9��l��m�Q<���L�1n�d��$�&7S�8Xێ*�/5#}�V��&J0e���HY1�{ K=N�����Z|KB���E�7��I��m��4�#���,�Kϻ\�GC��5�R+��QI���H򒚙��r���B���7GD�d/��˫�H��w&�q�|��P�+��9�/��q� ,����;u�P�`U�V�f��<���W=�[�Egl��2�$}�b%�5kx`T���x���v (���B�֣~�w1�#���Q�� (g��>��p5�2Eͳ!����|!�i\�:��N|E_-���������~:*˾�y7kgv�]̊���1�����9�[a���X�5���'��.��&�'��_������' ���|��f~Kb��J-"�E�e��oP6c�X�:["�����GuZf�Z�G�~���o��P� �}D���)����/V;:�A����w��9Hp@4	���/�8F%�P��-�r~�G³�y�uߖc�CC2daofEoE��G��C�`	t������~���2˔���eX)����]I�R��'yҁPH���#�#�����s������c(�d�s�9٩��C2�
H������z�#���y5���.�ר��j�o%��G)A�ৈ����r����v*d��Lk����v�x����o�7i�����������c��������4���l+�v�}�9�0\[!ҞC�~�;ׅ�ة/޺�w!��\�(��'�4I^G���0���h�<;���O��6�'�S�a��Y�K�vއ-�@�P��AohҐL�$Y�k>�He�w���3�}�80X�;'����",C
x�~�KrhЂe�'�.���F���l���!�<������(�w2�"�t�JB<��*�2J��(J����p�52S+���%�K�Ht*B�EV�mp�I�\�KTB;>x��L��Ș�<6飧��cB��7S��O�ʰ� �:&�����P3�����5F����S��ѯą(l�&:8�2��Y2�rB9B:E���)�S�%9�Z�eKD�C�Z\/XndEK#X�@T�V҄�[���ՏY;i��P�K�Ȱ-2� �M��͵D�40���1;Հ��e~�b[q.��4��TOl��LV��k�|>�NR����6<a	T��*o�R6���MWz�����4|�����8�G�\o/�𦵬R�5f_�͝���n(!������`� z�j����b��]�䏁�{��@�5Z��΅g���(ZH�U��`@�x�X��a�Q��c)���cENur��S� o�]�\� hQ���b+|�a4�:�y�i�o�-'�#;P��{H��ωk{�;�P�������j�'��;�(�.kq��1��#1� ����Ol��������#�d��U�(M�U�Q��z�M��><7	E�%*�E_(o��;�l�"���\gtb,M�k���������"��hV�z!F$��jy�jo|x�+�4����
�RS�*
�ǌ�Zz���dՃu�x>!gΧ(�~(6$���K�a�����41qO ��^�l��"���e����[>o�P�V�~����}ZP�?�A�«��O�;�A�]�M.�=>E��y�_G3��=9E}�V��Ռ�2�-�h��nG��*,]���(c�2�b}�0���W�"��BL0ʣ����`�-	���g���ªelh�x88���@�[k]�Ub�t̎�7Eu��,���em�W*�	���HX�Ad��q�Ъ�:r�����p�s" ȨJ�6fـ�irA�X��2���h�޴9|�SjIweBaD����
�Ye��u���g;^hs�I�e� ��Vh;)�����b
�[���J4��O�]O,BC�F��<3����v�4�[��p�8y������Sh�&v"sA��̆��,"��^���X˯R�F�L���3���Rv��5�t��<���Qpԝ�c�=��I%%��1qi?�����I����a� ����.!��,m�I��Ⲭ��Y��.|A�f��!�AK�-�v�Eq��G�>�����k��o,L�b+0�4�.,���.�A��=\�� ��R��b�%�û�Zm/�ķo��<�_���F�b�p�2_Qh3uc�wj��_u�x���dLL���&�z��z�t�|�-=�/�o�O5]���8l���|�ڏ�-�/ �bx����?�%��_�Ka0�i<*PMw��\�q�&n<��1���B@���lG���N�G��>->\G��y�:��x�]��Lژr�ye��7�߅���}�rٰ�i���G�̡^a��U[����/~����B�a=��;��>��܋`�/�q�{�yV^���T��.i��r����m[$Ht���,ExĤy`]/sO�\��h�X���v���q/��/��L�Sg~dߕߍT��9��;ˬ�q����=r^�m�	uAh=���)5�f�,���n}����Y�����P�w�B��>a,�:���Y���ޥ:�J����= 6��Q�DS�
S.PP�ɵ�4�J �ي�i�c���`�81�;�@�a���۸� ~5It�� �W�ڮ걸獋�	�(�g'���9c������ܙ;�v��t�O�?��Vlxf{@Kp�w麚a/ʛ�ZtD��&����ﱟ��q��5α�X~�&	h�����GߑM�f������ցR�̛|=H|E*�^��8�[��]_��4H\�������^�C`�"��t�9�=�v��RH�ZFI�mj9!�P�+��8�1O�<ݒ,�M�*I^l��;g
 fDK�j0P.��H�5���j�#��]�� 8�A>U*y�
ts�-"�6�؛[݋5C^�А�xA3�2��:$C�.�}(�i���s��d�Ł�.���&a.�e��_뛳eq���B�M�!��w��aWQ�$<�:k������k�f���]��hF��Dڂ���8�˞�-vbd�H�$�(_]}i��fuP����$�0�Tb�0��+��I�
���~I�V��u����	ޔ��؄m���Q�+��<����ݬ��� �P���7���R���d4ʫ"�E��!
ڸH�XwJ:���<���O�5����=��O��c�=*�v��e7���a�1�6���Up'�8��y �f���� �ع�	UU��~ӸI�� FW��R�8��W�N�աY���&�m��U�w�3��@��6}�Щ�]�[~Ғ�p�2>�c9ı/����v����m��KǺW��)��ᄎ�����F�T���?�yTT��K^��s�*�`1�>�\ۂd"��EY���!�oypue.e�e]u87,}�4� m���3�i�_�HD��Eز(��8�~Zf���t����K��O�%�d9��,� �=�
�:���]���1h��ȫ5��w%3�ciՀS/�AR+���3��2��� ��(��f����U'��8&��}2K�����oΐ�A-8��fk��_2����h�Af�/�rl���]�͔Є*��j����Z��A����9���7�p���i�x�8:܇ �cM���?־�#��۱�JQ����RKX~y��tٍԗ�K\YI��2�A$�M�Ϋp�-^S�{���~0ԥ����V������b���W�Nx��EJ����U'�r ��͌$�
ϻ�U��e��-�
0��P��;���&5-��ңáwdj�%��[�	m�?���g�����q���!��X���V+����x�V�3Ä���@E�.���|�1��a�]�(X��,�M+ojO�c��m�W&L3��w�x��,�a|W��×Q5q0H^���x]8�T�t�����l�Ψ��Lm�j)��4x�A��
( Z�7��t�� fq�\7�ϳ��g�H!��cH#�bs����k��6e&���j�c�۬��ґc�!(�7�yX���z+c�jE6&_R�7V54�0��W�X��VWv�ɻ��
a��1�z���|�1��C
;rL�p�jU�!r}영:-�^�#�K,7H�r���z�Q���	��5�EVk�>ls�Xp�u��g��Uǰc����&����03eL$b�������vGe�ŧ�Z)'
*���=K�,���+ղR���g��Dg�[͠�rG��^�G���xa�![x�����������F�)�_��R����DC����,�\���Ⱥ�&�#5~sY�:h�����H����$�=6XWtu��j�Ϻ��Z�uMJ��D��Y8(e's!\7�B��(�6�h�IȺ�����G(��}��+c����m߱�x�1
ŊM�v��B `���s:�b�{�U_��.��I��� ���0����W���H���m=�z���`r��̆��]���<{�s_����^ٓ���L�f
�]�������0$)�Gs�l�>�{V*��;��� ��q��Z@eg�����Hv��x��R��~�I���=�e�W��Q �U8lJ�a�to��BV�6��\wG�]�f~H~Or~�` ��Q��.i\�@��|	�J�ߙ�ni��5
���(=�m��ϯPG�z "����gH;�ռh��B��SW�L��s[�0�0���ȡ�~Isl���� �,w5~�u���LnrX����z���Ew�C����Xq!��{ҬÑ��".�էzt�+�,#� �L��b���>�Iħ��޳/F���V�7
�?���[�/i����5"��<��+�pC�s�S�"�{��̆�`�˯���bC1 z6������&��ʅ0I�[�4��umY�O����9�b$ى�WU9��c~g�KhY���ZM��*�o߷X_��ݲ"$R��kЈ~�*��XBY���Y�#�(y�	U��O�����#A���z=�>��$������3���,�9g�{ �-6Xe���̴F��3ZY ���Ot�����cb��Z��$�j
P��!�R�,0.ѮLFUc��#K����� ��q���K]�5���c.�����tqy�	0!S�CCZ;Qb(�i��LM����^���	��ѡ������p�8��m_f�ΰct����L,]-�7e��}'q�44b�{�%�[^���&��-��J�������uv:���'@�[��^���:1>q�5���L��ό P�o��#��T,�%�����{��N�Uo �֩|T�E.�_�C����+p�eE?�p���F��ɡ�jH�x�5�dVX��d;۶�J���InS0����(�(݌��k��ԛ����{�m�n>����eK�Wd�޹ �`s3�n��b��V�^U*���x~��{�[�h��ξBp��:�({���I�~�e�����n]�%F�-=�;�`<[��3^��r�?\�k/��
�0���3��� o-J�H�Y�q�~�,�[�������}{�0�h�+C�k8�t凐���xri�x���*y� �̢�<�0��ן<CyH�녝 �l~�-ٓ�Q�
w��4H���q¤��f3L^�Du���U�k�9�s��\�A��x� p�Tiw�3xgq��O�i�J�c{1��P,J�{\/��i�R�sO���*��Njz����������u�NpW��R��۹Gx��8�"ո�.�� �2��좷���ցԶ%ԛ��w�v[|X8o����t6Om9�yu`G�b��B�2�i��G#�3�1�A���$'��+����!|V��/J��~���SK�����ô�xF��h*�-�}ٖK�|X8�}��dg�F���&����B7r=����{�\����`�@j}��"8q
7�WHr�fˆF�	Yx�̊��X���pfqrZ�;��4�� >	i���M;C�w8��%G�ǘ�3�Ym�Ί�G�Q������P��uTU��/�l�+Zp��W(޹�	�-�%��op����Fv7�+xV���	�X.`3� GB��B�T0V��=Ѥ����bCW�.�W�r�oA��K��'Z��6�`�8!�ßx/�zQ�����c�L�'d@���_��5�'���$�N$f�\�P/�`_�#Aɳ0E?"b��Q��=SBU�=G�}���4 �Z���L7Y�������0du��|���m2��n�N�]�Ȫ�Kl\Z|�|���&GȨ���l&im�7�������C
caE��eZ���Ѥ*�������~%T�sKՆ���X�<(�4�����;�dH�n��3�vrĹ�冫zz(�Ƹ��G�k����1�>JDȻ�(+V��om����:"�JE,�=f۩+��с�:GgMñXa֢�t��L�`f��+�mm�V2�L�!.��=����纱3W�*��&5��j�_�����E8�f�mYl�(Z`���Kgi�7B���戤���,�n��L���J��mj�z�J��	�Ň��A^�('ٓ�̶�l/NM�bxcC�����,0C����vX� �D*�Ђ�,���Pg#���ūE�ǎḜ�R'v���:�+��׫m*�е$���S���K�M �=��x6>C_`^Q���vD^����n��Ь�,����T�p�{��ӂ�I�=~k�#d��wӟ�4'?�����}8�U���J�3<#P��r�W�7�xeuP��f�5�v݃��}r�*WA7ff��W�V�~R����V�
V-�s�0[p�.ϧu�Q؅�m���y��"7��H�gMCݬ��2	�+D���q�8g����UTo`�RgZ�}~�	��`=�ӗ��:���n��K:R|�bJ�g�����U���҂�o�)�]��`[ݍ�=����O"s&��� cwM$}�ORk��o*%�#��f��\��e0C�
 ��CWVc��v�)�I�h��ե~����d�^����E<;I��iy!�ߌ����J�����7l{j�H��g��^��w��]"l�Y�6�'�my�@LW��PI[��&=���?���(�E@��9 T�����|�#j��Kw90X��� �u�ƫ�����˽]���#�ߗ�9Ӭ���t�+9�B��D�I�Y�(��R��Ꞡ��V�s��J|ԉ�]�[���'�O�HBs�*�{�#��8 �GU,{~�����Cc6ϗ�Id�Z�y#�o����2��VyK�X`Va,��C\�9�٘����G���Ј�j��h�P+L�UQ�%��|7��m����{f	�]�� e���,h��+Em���ˬ#�s�q�B����3����y�b�K�^y��ʲ��[B�E�,�C��ⲟ"�}�I����]qG&uW�%�_�G�K!�v䞻W�P������7�]���}�z~��"������ T��7HY���^ڀ�g�ʄc"��iy���M��'��r^����,o�Y����ɋp�N�w��R�3�'j[օͿx]i�޲��R��6�<�i�$��K�_�w�j _�%z�Dʃ-@P�m|Zj�����bi��;Y���a���N.ҔX耗��B�s$��ˎ}W�Ӑ��R����1Ă�E bTV�l��[a�����iC�UXMt���p6�m��A��`*��(!u2Ά�z�tӯy�Cd|�n��9f��4Ԫ�YL���f�ٚyxa�%����+#�����<R�r�,i"�����w�R��U���D���ݢ�r����bpl�Xϲ��d���l[�ɾ��u�G@r΂�Floh^�k��l����y�\��m��}UK����`�y#p}�߇i���K���1�h��������!E�B�_ �6�= �#�c�������:I�GMA��"6��E���l��n�.���؁V����9�Z,e�y��n�ˮ�m`�i�`��{΁���&��/��i��:c_�͚ ��hU����E�۾]b�{��ݸSn�zA=�K��{E��Ô�()}�~�q����d�qaj��-V8���A�P����D�-��0ȸB+��SGBJ�t�<n����}$�&���h�Nӧ�?WiJ�{�Q��"��ٙl??����n���u? B�w��|��׆�����4�_�}���Am62q	�}*�2*��z���\��޼_�R�O&�{�L���ݼ[��H�b�o����rS� cP�[�Q֔%������MW��k���&{�H����th
�paHҎ��ܮ��~�����XI�@8&}�pUw(���lpb���˜_!Bɧ�J��fqP�����$Px��|Q��/����ϯ>GMı��3j�}c>�����������%g/<�V'���l�*�Xo�˥C���;��5)V�2c2`*r�g:�h���v���������@�����1Q��o���$�b	Q2��?�Og�b�9z�k'=��	dx21	���[U���C�}�=Ok���=��1�\` ��-�a�=���]��O1:�Zh���A���ʼ��9ҕ9���[*1�/�?��s�(��� ��V.�ICW�X\�G�t��]���<��t%s�Pd�~�n���1�4���*=	��z���3�Ш�"�\��*wt��)��#��?��D_�����B ����QX��ke�����c�ݿi���\������Q��c���j%��QQ�3ezȰw�Vi-Y`��çޙ��9A�{�E�=R2!v%��\+]�Ì�x}I�[$`�Pd���2��*~~�}�Q�Lb�-��1�Ƭ_F�V�AM[G)%#G�+�1��QylF� ��Owz�b�te��ޘ��22o`����ݚ��LވD��(���$��Nxt��%����ik��BAJmz�Lx��������H.�!�[ز�A)Q�����
�N�'�(��af��߶��$oJ�]?�s%��~`y�����f�2][#�FΌL���i �����F>�1�Ud�L> ���C���3��<�>I\9�Ly����W���@L�>�K��V�c��p'S�.�0���ӑ�0���h��Ѩ~(�K!_�$I���]7�7�)\Lbv�����aQ0�O�nn�j�\�������.=��z۲��Py�do\��h��%[��a�`T�ɒ���m�z��y�i��u|�2<fV������X#1���%�?5u����*��,�]v
�%���(����	�|�4�eY�?�*ڭ~�if�Cu�G�hj���It���h��<3�hC�{�<X��fa <��7!���Q˝�[K�B	��N�a~0йz-�K%����˳Y�axzJ��}�|�5���T5��n�M�����\�\���U��q867����F	x'/���P����-~�o%%�\W!u Uf�'Oٶ�����<�m�[�i}p�t��Y��AC$��P�rͰ�p��l��r��a��M�������-C��oc9\�%������O)�(Y�ٳa�bf��@�^�ꩼ"J�[��-���q>E���)�t� s;[R
�M�9}��EzaV��MD����!�a�7�@c4�D�v�k�_g���]�itFR��sV�R9Tjo�=���^�Zb�.�%���]=���ỵ��{K�"i- ����N��?��T�t��ȓ&��\��" �� X�P��[��VŪ�W�_c�g�[���.�����|�P7�?�C=��җg�˚HNihf���+��K[׶#%=��S������E=z��6c��R�	�ȕԿ�6�_�]���c�~6�����b�%I���:�^���9��\�>��y�7�Hj���O�L�e�xc�;uX!�r�)�M��V,���o��SC�LJҭ��"3A��17��N�Md���AT��t�%w�fW�B�{e�S�H��N�j�H��J�I�|���/d�R:\l�C��i�p)����h>�� �a�M�/-f����$�4��pY޲��#����{��F�x���i`W/�}��j����m�}f=�r��T2�U` D�P#u�m	���d�E�d�^zpa$�(3����Ş����?,�rI��˩q�i����[�OWV�^	�Ѕݏv����w�;�c��@E����׫X'D���E���)�q�.�e"n������@��˒�􏤧���ʚ{u,}U���	8����ѪD���������dP,�h��oN�b�\�,e::\j
�U�tI�-qg*п�Gᦱ !R��,��Jh���u�0�h?I�ܢ���=��l��>��w8K>�M�K�����]�k���ؒ!OZ�`�1
W�;�n��-D�z����;v4�����{�f�8h(5��͞O}s��t9*�3#�a��H8A�y�g��R1 ���`��r<���H�D:��Y��?���=��q<�7S/�m��������ڝlY'�
��W�\�_��#�"@s�o=���?�ƀm�b݁���t���7��L��N�+>oy�,{�!�Ƶ���m�l�!O�����9U�7�&����)n���� bM���(�?9o�Ƥ<z�T���������ˋme���B3O�䠾۹�i!� l�r��1�b��B���6��x��Z��qM��*w�� ��	��J��}�7�^�<~赚�˚2��~<MB�1u^3���>�*�^���3>R��lz���Ӯ��9�祍�ېv�UCZ�c-?���g���l\�G^I�>]�[?5�e�0���*�V�#��7X}>�̢��ߞ�e�ϓi$�y����O\3vH#�&dt���e��s��ԅ�W���W�\��lA�[m�θ��r+�_1Q�3L7$1R��8h�^k��L�����}R��8p��(Լ82"�B$����r��fC���,�2�j��� �i�˙Wd�X��2kW�'�E3�fa��&��u�,�m݂�� !7���'m�lY���%���D���H�瘀q"�e�x�\�=q��nwBb��Bй +Z(�{��+�W�������Mv�c�/5S�9�Dњ,Z� Je
5�<������I���S�@8%c��ā!z�̈́0�(�Jg(���|BPg���9�w�F�kC�6SA�N>�$��$���h����h��PS:��Kwj�]�t�C���� ��%�i�R�մ>��ͧ��?U�\ �}	��82��ǅ�ʢ���fQ�V��[����S*CStvY�|30bM�pd������t��woB�>��s����D�[S����8Qñ�-�&,rz1/�Ng���顡a����L����=Bj�H��t=��UE^��4_���M4"�����M~viw����?wy�iN��o~c�4I{a���uI: ��Ξ ,�E�2y�Ho /C��p都����\�Tk���vLct���:XL:�U��y+	������4+_�=���*���4f��:��fu��y�b��Q,p�k04�����x�g(ޡ������X�IE��[!Y!�tk�T�{��N+��|7���M��U*��q��[�������U��8P�P�bSg���<y�	��E(��sj�Vf#J�"�s��V��<�1y����@d��Z�ScW1���N��W����Ƅ2��cb��-_emUl`NT�l"�~�b�M�xiP�.�(t�]	��d��	�U�C$-�Q�yܿP���L�؜�5�lWEqA���\�����_��8mXySQ�z��s��z�҅�ŉ���yW�!��R�O<��"'�3��#AW�s��"�]˕r��{��U�OՆ���~H�tDM��rr��e�pMɱR�O�c�=�e�oh���)��!��]��I���'�Y���C�'�HD�@�-!�AL�ܞP<Ic�J������ʳuG��|���J�$*^�e�o�.n_怲d]g7�MA@�/>�.�x����v�E���cK�_�
�{ZJ���Y�q��q����#�_�E
���	�h�ړy�B��w^7ъ�*�栋�ٶy;�����=��{�z��/��^������k���)>�l�3���zS_�@0��_Ԧ�4J?�y����}�Nu����o<cO����Tl�#E%gw��	(����:[us;L�Ż?a�Kl�]����y����vIc�.w�*b�ҽ���<$s�OZ�5yy�x��6H4�EIw%��<��C��P��ӻ���I*�E���e/N��0| Ux�=�0/�U^�-#��h�;%uh�x3���r_�P5b�8��?�i��?CO��Bծ�L�ƍX���������8��s�^�;�w�D�����fl�r�uh=? ��OiyU�|X92�X���m�t��P�6~���.��oe���yBkw�"�A܀	��֒�G\�rZ��3m��3���)��%���fs?�ٯa�-��V�!1�S�� u��kz0���\z�Φ�8� r���Α�!m�^?+�^V|�r�%{/�қ3=��
��#�ϭ��~Sȑ
�	�Iψ�`����ud�ܾ�N�z�u��������Q���ܼJĳ�a����`�1�z�z\������s(�1����x����z}�$��������I|!@_�����L+Ӥ��c^N�
�Du?q)AG�4?����o��	�q��Y=��H�������O ������GF�Ce[���Jȏ�||�'�U�F_飚����F	!�{	e�Ɩ}��g�!����,ꏭ!}�e��kaT�.ފf��	���r]>�7WSW�|���>�6��nF�y�C:(f��wrT�k��\"��ݱ�V������*�_{�bf��b&�ԔnJ��Н���P��>�3��T�!�<�K�fy��=*��ř�4	֦g������A7&'�C~��I=b*�I�|�?��ʷw�u&=*���Y�s�}�~�v�%;e � ~�,Ob2A�6D��^�os�ծ6��,\u��.�E�c6���k\6����5grCPT�h�l+�Ͻ�8k�p>���^�4N�J+���*R�U'�V�ZtUU�;ݜ��k	��!�y�@��q�����M��WC�l@Cco�{�.� c���KPt/��UL{$&K%!G�I���L,C�z4��#�+L�'PT��	Y(
�2�:@~��n���猭~����/�0��h&����_
�`�`�y�;b��q�v�yu_f�Ay�3c Mc��h��L�x�H�����h�y|����Խ�@����%��`d
�m�>���> +�m'���|%&&��ݬI���&���˩~�0�`��,��'x��&v���z�/�[m ޣ�x:Dx,�7f-�I�(Xn���n6,+x�~X�,�}R?��9g�"��q�$��e�1�^�~:��|���<��d���)�z�/[!B�4vKLPڇh�Z��oj܌�=�R���E�!�"�Aq[��.��S/��jNߍ�nx�}�|����5�k��1t$�4AK�s<t�k�*�� �6�1�4�J�]��::���(=�Q�r�;��^Zt��bvGk,tk%�+�#w���W.��5� e���-�$��U����}��T�nd�B6��ğ�Ȅ�?5�������8r�N}��RT`�*v��<�X���~�H���oYh�M��������aQP�������ȏ�1��(/�ܭ��W����A����)Xi+������ؼ� �^�I�`�\^0��i��'b16)_st �tu�?��
�W�ڥ�g���_i0�˱毇ص��'� �[�az�9�}D=���Eå;pƬ��_x)^yѓJʷח��q�W��$X��Uג��7:�r:&-8"���^	�17�Y)Lԧ���M�� �������m���]�� b8sJ����DO߰����On"b�_�^�g� ݽ�[%I�ۯ��/�dD館�ՙZ
��>>�����T}�7&�<�;���J O�ţ���3�v>*~��.���L�<�qq#����iz.i�b�K?w��*۴���A ���L5q�N��!G^-@?-[4��C.���o��4���N�]X?�'���{�R�5���B?~��`��A�ᅏ7ꀦ;�v�^�r�P%� F���N/bi�-;F�xCg��� �k�y���K� ?=nX�d��$�œ4ݬ�w� An$\a�{��4�u%bA�i�!��L��8B5V���q?#�&��:��N�8�5�d�;���P?�OM�S9��ʖ'�՚:fӝ64�j-�Ğ�=ϿUjy�wΛm��z\گ��z�{S�7�ڲ�ऄ��6�F�M�j��.*-ո�gv�� 	2Д�Y�#��U�Z��VC�Wv*�u��Zr�|D�D,��+M���Vv=Y��*�oG�,wǦq����^2��B���;r!�Nq(۲����p�6�,8NB"���o��؈��P4�9��x9B�܉�:e���o5�����԰'�n�h7����<Z�Ġrގe�r|���ô)��M"cd�bez����4���@�D�:��7�I��{�#5� 4@�~l����0rim�acW���Jre��*�'9W_r
��X  3x�B�[�?�7�yҗ�\a~_��yO�8t'�6�)�?'硠/�1?���}$
x%�Ü�b��';�AR>�� ܮv��p,L��� W�76�R�6Eޮ� g�c�"o����\Ă+�r��%�m��,s��)��i"6[���w�0}������d�Ĉ�u�Py��T�|+���/�^�ב�rzj��O����S�ߛ�ٰ���I�/j!�w8�.o�������y%ĳ2nM�;Da�����}�bv�<36�����¯%_p�������g�; nQ�9?Z�" �ê�g��־:,ʔq_4�)����ti�k�Ӛj%B"%!�C�~���u�a���vΖ��%�cnrH��2��8I�?�I��_D=�x4��b�n�q�p)��x%gn���iy{�6�U ,��3%O�ΊYh���(�m�~l�Lg�g�5*�@?~���P�����������~��L�ӆJz����g�r�7�I> Y*W*�}�p�P��x~&޳�*�2��*�+�$j��XժW3z���-������Df��w��u2��~��z�*l�ѓ}����7D���r�=1^|	{�%q�7�Z_mi��i^cK쩳�HM�[��\�M���ad�$_��%͊ٽ���O �@�9�5/��Y?�u$t'.([�X� )��rw���Ƈ���-L�[�t�~��&8�S5���R|�*���c�_~<�.E��z,#V �O�e{��/+>�L��R�F|/��7[+�?xu���4�������.�$���0U��#r��Ø[�s���<��T�����U+�����w�Ȕ�"FΕ�[�c��$)b�I�n�-���<#,%�΍A6���������e�zO��d�N/˜�4���g���鴹��:���O���~+\�
��W(.���!����p�t�qs��vhC�4Dřurc~�l�&�6���=#D�|9J���t�0�H���5��K\�˔ r:Y��CL�ww+����o: �H#��nA�壆[�����������, %�E/ϧ�?�yM3/���L��B���^V:d����Đȿ��@jl���لT��{T����Z���� ���b�̨#^Gk�,(}�N��w	�[7(��û�{��]0����z�]���y�)K���e�B�*�&)�9'J4=	���h�a��k��4�Or�R6�.�| ����1�],e�M��^��ߍ?M/�R�Gi��K��TK��Wjo=��m�_*���^�0�_@g�ց�0G~�}u�@zU/W��&q`��ym���RP����8�q8Y� Y"������3G�G�����+u�#�(i]мC2h6�5�ʺS�L��+Y���Ռ�u~�Z���6�^^�M�<��zR/Վ4ݱ ����J������.�i�-%w}��'���B��ɝ����o�T%������_i�0ko{@D�|�鈸E�}��=�M�Y�L�_9�X���}s�Lb���̌I�
�F����]�KO��@(}%�H-�3�E?�v}qd�����K$�.H�h+}nf5�$����=e7^�-�ޮ�ߴ��&[_��}�*J�Bwi����� ��K�hC���L��6�.T�<|�Bbʎ�#x�����zv����9ʊ
_T��W?5Db�	�z����OO�u��('�$�&��6u����I�Rҕ���:�J�3����k�ruc:i�@����`�ysi��,�!��UA�V]�0�B:҄���!��	�X���C�(�'�@�ܢ�kq0��Eo�3������,�7Z����OOAe;���޸#�\N����G�������9�$L�����qb1azc��y�t�F���o_�P��RXڵEsx�V\vBWȜ�` Z'%6(�;Z���U/+��]�{
��IW*Q��,��)�l��Ct�����3lU�1�y�ӓ�m�w���Lm&�A�"�=������G,2������4~��HX�)��ȓ�2:�q�#�H�`��i��z�N�ʻ��H~��ߗ	��w�����-��I��m��I ������de��Ex�NW'�N�`)��ެ��F�ua
n����v�u`}EO���t5]�~C3�����c�pZ�"�e%4�l��	*jbG���S�g�zS����W�I�/)���6�Vu�bd����]����;.y`V�ݮ^���ct#	E�{e��9��A޻� �:l�ړI{I)��#����9Q(��f��_P�M1lio�C���,׈X�s�J�)d��6��p�2���wבj`3�1 ���(��8t��{Rx��$�7�4	H6.�f�P�yFF�q[��wg%�'�����.h~�=}G���h=M2�.sLޣ����<�	>��*8/]�ڵ����Y�5ڙ�01�a	���1xqq;����@���c���	���*�l*Q.Ժ�haG�0R�ԃ�^�~�$8I���W��t��̻Y	Jr��1���#j:��%i��o��x��.QC�%%xB���G�������]o�D���vK�]X5��9%4�����C�L�R�YňLJS���#h�U�EIJ��h���0w?�P�?��o�`�\��{�߮6�62��,�{k�s5<A�!����+�+4T��U��FOa��<ϝj"��|4<2(M��;��� ���o�g�(t��1�j**�1Sl}�p�6��a��Z���xX������$p� �����a6N	y�s�-:��Ct�O	:�z:h p���W�����qp ����>N�9��.{�FNa!�hVG�̿��*X�u�\�h�����9�NE`K+W�{��`�MT�u>�_��i�<]bKY�X�����_{�	�~�V�'�U̓�g ĵ������S�M����3���81!��T��	�f���4�������Wk���5C�[��D� 'ϐ)/�|H�����y��7~��f�΃�u<m���'�M��B)*����f����YN�=�����Р��o I9*3��>i�4�)����H��j���	� �{Ԅ�ih����>UJ�n�&�؄��E�)�j� �yܚ6�)�s��!�3ւ��"�����Ȇ�_��>��٣��I�(ν,���\�d���sG��0�����k3� ��� 8��V�_<&�Yk�HE��Um-�ʹɪԏ��3\�\W���X�vo<���8xaV�sb��l�atA:�k��������̈3��Wd!^�$�Q�qois�>��s]p�hh��Ǎ~r�����g��1�t��n�k�:�DF��8������y�l�ͅ����w||r�|�^d#��K7]<ΒĖٺ���ך�ya� R|Pc'p�r�`� ����f�G�1&dc-s���d�Ou]��Y�Od���7� ��GN-�B_$������@��RBfRڵ��|��N2Ċ K����MكW8�Ob��键�o��A�u	@8n��������؉�����?�ov�dX�`���������z�e�B>�_�F���{Y?It�U��Eس�U �i�b�}H*�X���O!lO�UQ�6�Ǫ�8ײs����0�|R2+=�_�4�VM����nUX��b���k�Mk#;rR-|��AT�}Bl��$V�}s$k�Y���W����ⴿ��I,�p�Q��5~pV�'�@�'��>�B|�R�q���]n�S	i9jk�T����k��ד�k��7"�r�3��p\�fB�xm���]=D��3U�[*_`	7�]Ct�)����9��*2DōW|�J���ut]�:���^��U��4��H��������G7)
�v{�J(%	B��x�V&9�����m���ez�K:��iX�'{�'��[J��'��/�S�C5�� �w_�) ֦:��pϛ~���@��\<����֧x��P$�3���u���'�>/u<+X��&�#�P�g�wZV���w�{���cfۨ�L�[�&��P�[�I4�p�ͪM�c.��D�+��~*]�6�޽�U�ߛ&�6�X��9����}����ҽ��.MD)�0t��Ϻ��q��s��6�=���f��W�1�=;�|�#ϰ꘬���	�	�8:J0���W<��2l�+\��=��	yZje�u�K�%F�6���gy��@��S������˟�eQp����T���Tph�g>,��^.���Fx����+�c���~�sRAa�����X��8������
ZB����M_��lxd ��
,��!{���ɯ�'x��x?�iT�Z,3�>�1K���L)2~�(�0o���%.���	+%�k�a�@�^�/
���4��;�b��w��o	PM�E�&|d�G��<쇧99������P05�����j�<=]��8��(J�%,!�FJ�6�ê�-S{�G���U�S:,�#�����o���g|�s(��v��m�횭J�gJ@��?A|�ФSԁ���!:�����SU��*�^�Ԕ[
t�"�.��1{K��$����P�>A^��4��lLl�5h琘�<~�1��y,�q�q���rLB[ȑ5�4�n?�:�S�S~D]{� �{��5ܭ����T�,���t�M�ɇ�r$3��U���M#?p�ռl8̌��^Dev����Py�^h�e�٠N�);��*��O��R�Ak��r�h"�Ϟ��7��Q��կ��vO<���"\i�m�����ZP����5ˇ�}|��|CR� ��4D�S�-
%�b�O���՚��J�³������!Ras����-a�55�$}wc ���t�� �]�S-صH6���1��:�~j�@����3��)6��G(	�� +OEj�'/�d�>�uC$�J�����!�*�\�*dI̘p7wXP/><��e,J<Z:j���0ޢD��T���;RF)���2Y�!��t���kn6l��D�R���b�L�L���X����#�M+|H0��CW4�}O�q���&�K)�E��uȧ6��G�1vkQ�˰����6��Z�h;KxҒU�1���Q��&f�u�&$�D�&wQ[�o�u�ϏvfsU�A0'U(;-I}�����h�P̶��O�&r��bc�>ەu��A3��#;�x�{����kMx#�>�:%mL��C?�&���z�P�'d y3��b���8�����Dǻ�2䦥��+^5�q�*QP5�Huv�y��iҶ��!&�7���n
���#��UfN�o��� �`�.[��V�(�ǎ��&��B> }6�����8������9-�,��IF���Lt�FX�C����0[�7�c�7<:����_h�0�a������cfƹ=�I�GWyx���ǋX�k<�+Y����Ee�&M�Pdf/��o�u g�Y���^��	�x�{��,�o����GC?h����}��݅�.Avr>䃊`m]�]e:c��"�ë!��΋����L��=fiNΙ���c��J9�F�ND3:��"~�&R�����r���"jS� ��җ�����ܛf�l���`p�fu��C&F=z��x�YJ��i����%b����2�FA��G ���)�
䆶З�2��B����@�{����qa�>c� �P3#tq'�0J�9e[I`@�ʪv��zL�����!ׯ_ �`Բ�i�#�?N��M�`�)=ft}G}�Y���n��=\�ד�*����7s��r&q�]��9�.r�
��B�Q�ظ����˕L��4�A�6��=�6ڂ�)@kn�h�Gi��9�G��3�W�~F��z3���6$�� �_-w�C)m�;}�-2�%|\2����R��^-$[]�TÌG�::R�`fi���<8\M���)DY�����s�qq���8�'D��&�����rbdks��r�/L�m}Ԍ���׾�(-c��v����N������ $�mV��i�C����H�3���=�D�^5d���w"��
��-�眥/�8�3"�[��t��G���U��]�aH�Q�/�6�ʓ��ơX��W�����n�o���ң�S&��x���Z��#L��Qn�I\��@3��Ơ02�Z�Y�z�1��Q�Y:tg�v�)s�I}t�r�I.uK<X�,��(�h�l1�#�K�����Y�^��N��Lʓ]&vSǖM����{��q��Xin^�%44>F���\�YO�ϧ9��&�w�� �1'��,NJ�)���~�w�19Wq{��6�դ�z_�.p~�uehk'���Q_ՙ(	R΁d�
#w�L8�R�pTЋ3�-�"��Nɤ Ҁ��qs��7��L����%jg�23;�~~Y�ԏ�+��O�E�5���pn���[��K�hc�ѦD0>�M�̏/�Bn�6v��R�]3�����l�ϺI�UG�G�� ��*(��a�u܇le�Ͽf��2�0{���Mv�fV�=�,��b�9��4�i�K~���GU�Gl��MqԘṼ!�cpY.��������nSp� �~�gH%�1��U{�j�/�Kˠa3��a���Ō�G�Vŉ8��,U߼���2���K?��P��F<��)�\2�R����q�v���h���t�n4K>Ih�z�yQ�H��1�BH!:s�7b�%TI�í,�D�n����e�u8��v�OIC6���y��J�';��`��2E���A���"�8��ec��Y��m�\�߯��d��	�V�U����\�]J�3Ϳ;w�����?ϓ�㯺����]����%`���F�'���*E� X�_p~��9j���4
ڍ��3�%���o��#���u��6��4!�B�Gt�O��1W�Zpc4�Ƈt���}���\���Zp�*I�n�)!��sL���>�j	��twy�|},g*���]���c�]�`?�#��Y����W�T�8a�jj��T�F�F��b�ݑ��=��$�Ә#�w���n)^L� 2�=�v�2\If�������(#����w�{��.��7C������������! )�,o�%F0�:�{�i�	��o���Z�T��L+���ȗ�2(���ؒ��ѽ�:�t�h��纏s�K�lz�vB������,�Ρ�m|3��0��Ib��2��IJ�O��@~����YP��^���fѵ����������y��<����?�nں�Ԗn���j�CR�	����i�3�gi0h��p����D�^X(�;���6�5��=O	��£�s�*�Ƌ�I�t���"
ΊI�7�Y�6�t���H�d�
�Q�ŷ?N���2���~Y�}�Εvbg�(�
-ͪ�WzW[6�v����J�
�::#x�C��O���a���������T@!���ӑ�Ń�l��XU���|���
��J��G�S�{S�^�>��h�w����!�hn���ڄ7;��(��4�7�����/m�dP����A\�^w*�U�Dhxy��{VS��ʢK�?�^��~��rW���-|�)�P�((��HQ}x���B�� ��2#� 6��'a�q%v$�t�?�@G���L�Uu�6�"������Y�鐬QGyf�����+��g����_�n�}����⒖҅z�F�#:>=�Ba�T�OP�/.w9�p4�>�IT�J��qd��Qé&L���W��o�0ғ0�y��p� �I�y��6��� P��K��~�p�l��إl ��Yq=��x�&��*B����2�u��P�.�*���O��d��i�/����vQ $��j4@�c�̯6���V���[.j_ڤ�g�%?��_}��`�?�5����ڒ> �j��T���/,�%T��*T�GId�1�(Q~�6��D�ρW���������P��	�b)���է��`4�)6K5��!S�^rn1p�k�ۡ�Y��"a�;�3�PxFo�V��*Y�4%\��
�ú�b��i�H�5S�ƽ�;��Dm��5n��=37�0��I$w��PE ���g� 34��䴗���V�xD ��k��iH���/NJ�}�P3f�KVO���L��4o�f��WG(o���mɻY�*�m�;����
�HS�0��#�f�V8.�2i_ yŪ�ql/"��.�O��|�8��;)��.p	���!�@��A]_�eZu�UA �����;������zvEn��:�G,>�ن���J>���Z󗩄N\�����p��}����L�:�B�i�x�e�m�:� 8�c([/rn(������0��yx64m(`r��H~=���Pܖ{H��p�����>�}����XM�ѪD�w NԘ�w6
���v��F��,c��t�b\�S����!\o݉\햃ǧ# 6����/��U��@F<4H�>�-�F��R{L��LP���Zh��]�Ï��(ŗ�3�?�7��쾇��E�Ú�9t�W	�?�QC�jCrK�/&=�#EZ��*�m]?h�˷:��ι�IމG�{�]G�����N��79�7�4R-w�S��̑��5�	�o�(�C�\"��C���������B���j��`ӥE����B����f
�tE.�hSN���G�Y�b�r�W�A[cQ.�S2e�b�&��b;�/J�^��˜u���A��"�Ј�j0PJ�����[��=��R�g�hX���%c�+נ����u:�g?	�٧�?�Ξ�hN���_f�Ƴ�+����-A�l#�8�^�(�-���{A�G@e��a+�~�p�<�D��&ۋ����i�43{vœ���0�jۓh����z�$��vٷ�C6�@�d���R�����;w[�6�Ŭ5��*&d��I7/,ǖ���J�4�6�6��I<`�x�%mW;Mg�UAr��Ί^󟸜�xܪPip��|��9�}�=����� G?�ܽ��M����}��1ێtX����ʘ�9�	$!(CLy$�܊T�b�Y ��$;��	�t���BK�k��+D���T�pLiPVB$��.D����05��	����=j����M%2x�;6��n��Zg�&d9��kxl� ���yOjy8��ٜ[O���<�Q~�;F���T�OX���Q���U�f�^���E��^�S��d�G���7�S	v�)��?~uD�����:��6�$fa�φ�����1�o�8�;����=0� }X��a��Q��:d;a�̖_�����5X'���-`R)?oE��uy)H�oϏ�Cb��$���.�.�{O4�<�G�U��C���%�����g:]k�gI3�� Y�z���N=K� ��AC��6��l$��_�L��{�h�N 8ʦ�0˓�"�:߸p1['l[��-)1�-BA���7L�Q��8k]QA���vh��&��K�A]��]��"x�"թ�'�RO 4`��2��e�&����A��孟�>LΆ���9%��<	�=�{s�!�C��ԨG%�$5�jpx}�[��>j*B:A��}�col<N\��/��\}��x&�6�!����\Q=.�:��Dc1���Aݨz[��s+�(�MV�P�Fn#�
O�M�!��zV7t}�F&(SS�]�M!���Vx��Eı͊����쑸�����6t����l7R\��%��0�2��67z��L�һ䅥N��w���[~��7��-T��οT��3�������_#�;=��S_�	vp{��Z$����x�5�no������ʠt��� ��:x��I�&�L'`d��]�������}��j�i��LJ]�.���Md��vSUۿ}̩ƻ}o��h@�����8����0��o�驔u� �4���k&����,pz�tbe>�ʾ����ƐU�oi�;��f�v��1��p�p�!+r�G��=~���F��΅��iKh��0��Ԑ�钅��PT����䖩�Zcy��q켲ɹɀ��A�_�M6,Ki� �Նu�j:I4�+��hs^�դ��
su�&t#0�X{���@${�S$��Ʉ܌��9�O�$�f�>,t׳�������<"+�`&�NQ�Y�nb���~�K�?��ru�O��82��#K��X'S>}���%;b���k2��zh�vؚ�����������^>����C&N5п�ĕ�C�e7����'����� �L�"��)�9)�������������ϺZ���
1�ۉS�����_�;R�47˶c���x/,�+o9��/���,�pe>��%Z�AJ�p3ٛ�z�^�)��Q�];[��	���}!a+p1�3��i��پ������6�{OΚ�CO����5ߨ �����牏8�fj�z�yR��xb�� �z͂��?vq{!k��v���vW�F�l~���D�	0O�b�H����W��j�(<Zר;<�H�����Gs�b�z��� ��~�U�y+$Ԣ���$�6y�z�ΐ XǕ��U�Q�
��6����sQ�E5"Ct�Mc����Q6��	%�������� ��Xv5����raX�d��ϟ���%��U����.#h��Ȩ��S�w��n$�(m�P��0��W�~:[�8kFl��f0��i��T������ƬĿ�$�Hٜ ez.�N���ܪ}T#Ԏ�Ǘ?��Q1HqC!t�J?ȶ�e����+�$n(�?@�hL��P"�Zv���@35�/%=M�4Փ��ע^����'�)TCp�vt��x��s'���8���H�q�Lr�>��˙��u�<�k �V���ɣ�.�n�n2:�6�^L���D�#�ZN���!h 
B� ��-�w�9}x���D���)l� K�?1<��-���
rvO��p7c���l��`h���}�T<˻g+7Fi
qx��c�W\+rHsv$F[�Du�֘�[���jR�%�7��7��o��-H#��m��ɶ�sY��de���w�^U�].	O�6����D��ISM��l<�l�BvU��zL�W��"�h}��E�<���;tj��y��K�p���Ťdc�ّ��raڨ�g(�)�pZ&y�s�@�	O}P�m��і�xwyc�(S�g+�
+�eޡ�Rqe?��Z�8��7[·*r���vB�����h��E���M<�J��s`�rm�PP��D �K���< +��1�Ŵ$��m����J���<M�p������s��77�T��n'~����)k_� h~z8���Q�~2Tx���@@ԨI�9#4���~[�G�U� ��QHbd���%.�R��6�V�v���h�\�7�z�\�<}[� Nr���Cd�]_O��}�S�T�	��5w�?"S�ӄ��b�������t$�Ě��H���e��Q7��J��d�*��%#O�1V�%n�'����5��*pzm�Ϫ�����P����D��W�h�_h�ZCSr� �܄O�q��%� h��|�O�>��ϣ��N�	6�o�5=V_yr�B^Zv	�nrBE3ׅ�C�K��c{�'9ZC(
��0:}ӝ�~9)�~&}�3���A��P�_)��Q�d%��^���_�D��0Ӳw����9���j�_S��&�x��j�W��,2���ļIF��>��,\N8���QyuL�͗�i��
�r��6�ԥ7����ĝe+�`�9��P�W�1�x1o�D���U<ϐ�uז
(�f?
��&'�kN��?�����'�*u.�!Q�&P�f7!\�Ĩ�{�5Fo�q]8Ɣ���aZ���'��tH�`�� h6���y��r
��H�~R�2r��/>ޓ���Œ.���Xk�8���%�W9�vj���$��b��Ju� �[`#)VMS6�Qq���f��]%�W$��pJ�A�76����a��ss����5�r�b
o��v��1���p"?���-��5]��>���1;��%��	�Y!+�D���ot&����ҳy����SS�o�� �d7I��fx/Gz��F���o~̯�zN��;�i�C��\��T���z[A�o��df��S�L&Em1���F�#�u���G�Z͖榌����螀gx ���B�:\�Z�=��(��M�c�X�К�Z\S�ӄ����'oA��!(4����y.�o� �� ��t��e�:c?��^��cs|�4a0�$���x�{��>�U�P�� �}��C�e�.QW?��#��Ŏ�i�Y��AF���μ�Y���c_�S/�r=���!��q�}�-B��jA��3K�V0�P�FҠ�G�v�l��AQz~�ϠQ��[ƯUk����#�Y��@�L������:xw�pI�	��}Y�� [фZ@7�fx�&����)W��8���(EE���-����c-��"�F�N��f��L}s�ఐ�\wI�H}�+��h=X��nSN)����`�kO���Dr��u���U���lʓ�`M[��W�4ʐ��M�o9z��������[^
5 \eN{s�|�F$��)��-�j�e��E�Ҍ7G#��K�S:��Ik�Z*�`!+����>�8�ڵ=<�}����I] $�����e9*��]�Ff�)���z��SSȊ�%�0}�Pfh'�0T z輞�~�50�b0/&��o�Or�NC��ev��V{��{�
��K�OCl��N�kHZ�D�|k��ݙ�)����~��t�:���]j�c�Y�޳�1��"�u����&�->�Fg��(�'���l̜1�=���-�IN&8��D3�����1�@���!}�j�s0��4W �c
 8�N�L��F��}��c����0�tc���g&ǳ�UUr�-9��n��z�����8�7�]���}Ku�K�N}�:�4��Bm;ڧ�����+�-�����̅�f"!���w��%�B�Ys�5�t�`��mR:���TӺ9�:�`�S�dn�-�b��J�>��j�&��6H5�$3�Ci���؏{P�|���
�q.M�����$tJ!e���0ai�μ�A�u�[��	�[% �(�Yc� ���%�.z-���,�3D�ˠ��l��*(r^-�E�6alPi��2�����F
`���̔7���{7��Ab4���Iꖑ�E�<����E�Y�Y���$g���`&����A
���X�����X��_ln��_qZm�됗cTT"i��A"�͕W3�E@}��ʷuy������<�'��2)(��ʊRNu�a?)�����淫�f�K��\��e�5+EI���;��c��)���2+l���_��| %AA�a"�ݱ�M�� ��>�A��'b�� $.l
g�?3���?ě�G��B!��Ub$N;n3(I�(^ɷk!t�kk�~ii����h���LU؍Π��k��~A��Bc�S��BE��a'Q8Nj��	3�9�O�d����6H	uxZ�ګF�8�j� F��m^/:[*?���kk�:��)�J}fݺ�RH���(�|���$�B��ZB��sۚl��D�kY��9�܆6�;�t_�@a"�8�
N�� ��+�����sZ�gf���ɟ��I4�sumR�K��'ݖ���+ۋ�7��E�+�U��X��	!��Կ���}�3'���|K���J<d�n���-��(T؝\��F;*_@���g�\,:$����S4&X�)�5s\N�H~tV�䱢D��+�M����� ���+!ܸE���s7G�� �uri9��˩�)A�����L�������	)�U�T>�	4 (d�Yҁ���:j��hw}��2����"�׺ڶښMpB��D04��A�`��f����{�Ъ�%Y��*��m�Q�ɯ#"NO0�L�&�h��ݯ�����Sm]t�`�)��p���v��b�`�;�.��s�BR'��������h�H����h�SY��w�P��B=~� ��uo**�?!���O$�$�Xt��*F8�!-I�z�&��+��	�YJ]��`<��̼�u���`��@k�m�F�>�X���؀��.�b���ɲ�x�y�Hc���beJ�_����n�S~��aՃ/�q��b{5��a�cE�bN��B��� ����L;
���+!K~�0���U����F��r�q8[�Q&_��h�6�f�۞�_.��s����dy}J�~�8~4mRw�d���zx���5��@����Q�p�#�xO MZ:�R	fm�42�� ��&@�w��;k
2������+om�f!/�)~|�A
��n/��*-��SB�A�n�ء�c2���;�V�
@�]��G�����ߞ�LB����ƿ��h#�w��ED�6�Ũ7W%������<V�J��LK&'�n0DoS@CoM��{:�⴮��	2����dn���N*�iD�j~��ˍ�����̊����Nv1i�R�a�J~���޹�,Ru�W�7,عOL���>�������_��!0r�&�e ��V�)[ ���SW��r@)9�{ �e%-7�(��hCtb�*�Mj>�t�Q-!�{q�%E	���HM��hT_zd�д2�׳�V�޿>z�P(���HJ���@ǽ�
����˱��-��[�WJg_�J��&�w��g�t��]�K����c�e�|��*�9���:²�-����sK7$z��;��G���T���h\w���(����2���6{(^�ZL��8!0A/$�=����������<����W]ws;TxM�� `��cg�����>o$%/}��$��汋�jl/K�W٥�8�c��v���O�>��ܥ��m��:�+��8a� '�F�� Hw�_�Me�]5�Y�a�]V���W0�܂�%G�=zqWfg �Y	��#;�<�VH���
��`���e�M8�8'=�f��A��%��
({iӽ�Ykϸd�3N� +��p��W0:M$s���U3��d\���/	j��p��/�c�(S�r����K�\v_��¾v ��5$?�RళB�dJT�L̘t�����3�d[O��~��*�·�{���A`
h�q���b����2e�f%m��\I�=��T���l ��j��	t�(���;'%`%z�Ƀ���%�z�Gl�	 �(c*'��Zz]l_Ծ��?����o�%��z�Q������`�G^���U��OW�?U簾�d�#QtX�$������nk�	�F�������"����*,�g�B��|��� ��bw����B<��*&���^���xC6��b�k�����%�*��k;&e^}Z�,���#�	:2�he�۠���>\db�!*J�n���:x32h���E���>୧�ˉ�T	�?���S�����1�7fmj�z�[UO�c�!�(Oa��嶿�}��l�4��%}�8�%�50ǲ�&�f
b���d�i��ɺ2����W~�yy8L�S±���\2����,��Vc��[�+�Ĝ�f�	�XvT"���wsQZ�+g?�,r�&n�ܰ{�~,2k>�(b�O�� ?���� �X��Y�֘��)>e�#��F��[���p�J�al<�"�U��)+o�|��ǫ�J��@��t�D��wg�uп�7�%Nr*Ȧ����?�I�
����k�&T�r?�U�)b�%<aN�����u0+�fLn�����60�+�V����q*/gz�p׾�]7�����L���G��;n�`�"'���4����ղd�����'���z���[�����O�ɚ��uW�jh�g��w���:��������l^�k��kr�B;��\կ��MǉV1! �p��nД�4g)�[_~Z_!@��˽_�Ag��.��Ҩ�j�p�n�ge�I^L�#J�aX�H"��o��n}�!$Gہ�F��v�zVw�$����RJ_F,�{�S�����';�dS��^±P�!o4�"��S�Kv1��l<�����S}�k����M��'��r�W�aŰ���NE��G��s-�W;�zW�c�����|�Y��e�"銠��B��:��4G@L��;"�Z�3�[�+�Hm����<�b�1-�t�pX���D���!B�mm9���z|;��:r�vTa�l�������%Ue����Ol4�(�դm"r�dv�j|~=�W�� =@�/�\�S.I������[ #*�]�{y�೏9�]:��Fm�S��G�E�Y,K[T����9WI�{C��J�'-9'p�cͻ۞n���-e��gp@x^�;��*�Ajn��r��4M$a�'�;w	���-�>��J�dT��x�"dJ��A�f$x��oZ]"�ȎBf6�p����v�`��g@�w �r^���U��ߏL[�_��ѧ���K�-�;�`�M����
=��hk�ۓ���h�I�p�)*X�M��N��N�%a)4g�y�&����c�)�Y�UT��I��(����e�$(���tc1��'���T���I���en�-"�I����Ps��t��:#�����l�L>i�@��"S&���O���fsT�6����є���f�u�"ʣF4X��I�$����3=��Φl�-�̈�wܘ�;y�v��	J�в�jl#j(�=���K<�;�π97��Z]!A�o:!@r���h�wq�~��]�k`)��gIfk43o�Alf�����J���uE��VP?]\t���Cnj���c�=Tʑ�!�2ŀR7�M�Z�w����t~�)�,]��[{R�N�#0�D�m�>��㡓��Xϊ������{b���V����1c% hc�t/
Jg݉G5��Q�C<��]�7��f�텔�X�"V��$tz%���b
q9��Ie7_�V��LTk0G�lA%�^	r��:�@�@<���Ɖ�mP�e���-�z�)]�W'A=�=�-����M�yaZ,&�C�[�d��16ҷ��+b!�A��q�E��dE�IMxj�� ��
;B��ռ0Fx���d�}����kB�Ś] UD0�Y��P���ȍm��Fz}�b˥��r��b��iI/pA���W��u�hM��n__�ejs4m���T���چ�^^\����
�J��HKa͏�������A�@���$��z�A���(���
��2�=�nk6SO���#$'5��2~��I�*������w�W����ZI!�P�T�}�k��<�,I�׊s�7cΟy��<�d�U#*��M�,���@k��rd �!�����F�-�����ڤV`�T�e�^�5 ~j�t�}�7�D]ڹ��L�nzѽs�� �6�3��}v}�n�,K���|ܻ>�y���J�TTК\P�	����]���ݎ�;��~)Tz��Ǹg ƼH7D[ᯨ�B9^�Xƕ�Cw���<����]!��!6T�b�Xk�0�N��d�σKb������bT�z��@��υ��>�jŮ�kX�a�bz�V�]���̫�$Rͱ�$g�þK2�)h�@qA�x�9u��ETET��z�&�}#ܝ�\��)�����,	sK]�>�[~��}@[±���N����ӆ �;{
|����|�P*?��T����R}�~�hKBnS�2U���nT9OWVO��g��X~��dȈy�D��G�!���_��SGki}JQٽ��[WPkȷ�U�
-ڰ$%(Y���Y�1��LC���1��	�1�3��	�:�T���!"Al�Qt�%y,]^e.u�@g���Ŭ�݅��$e�m�I�ɕ/&�4W$.���/��K~�W<��z1���O��bW�+,^:yĸ4�:�hT*I4�u&ҏN���0A�!_���#�m��.��]��Z'B�I�C&y�)C�0�+콷��
���;���Rr�5a]��.���͛R�e&���C��!���lP�3Q(���0�L��d�:��Ե��$��w���_�>�
[vŇ�D��z5vp�	�KК��H[1?+����B��;���;M���D�x��=SrP�uI�@k�Q�}PT +BJ�E�-���9Yl���\��DP�jd���d���p�a5+�p�Ka��#�Op�;k�Il,z+30��� �����.@�u��;?�F���]D���w#n�{�ͼ���䬯�cJ�Ց��I�Vx�EGӀ��ypW��0��-�X����9
��r�|��L�=�-ZA�x"��ӎh�(�~ʟ{���
�1��с +π����rX*@�A��Q6#�T/���0�����d?���CE@Q�~��!�T�2�BD��h���V-E,-���!��9Z�o���m��	1?�0���L�؋���?z�K��7Y%C��a��!	�N	�񷫌�q�ߓ��;-Xr���*a})������ ڏ�4����f(e�|��5�Qj��~���L֑�Z��z��hЅ��kk]w�;{�]J8�ӿ+nǾ*�E�P��˯��]"�5Rt��������d��=�qN�d�f��L�zk���S݋�ȫ��#7Y��o�e���.P�� @���ʲ�L%��y<ZRg	����8�!b0N���O�H#�5�0���S@Z��#=nȋ\��B׃"�{(�k)����m�i�~�*���9�k�T�5+��-���*7�@�4��A�z!�@�DW ���;��lb���6U�\ߺ�L�m{��ssF#�V@����C;�UQ�K������Q��/����y���y�w&#,y���V�kF�Ꞝ��feot!<�O�: (e�� �-Q��}��J����8�=y���uyp�u!op� (����K:^��=��~��x�a][� 4HP���	������اd������@X1!?������B���~����]?���T߭'�754���p,I��P`�Ҟ<�P#���_\�|y�⯰����D��;�a����{d@�OT�������V��c J>�_��a[F��i�A����P^��M�_�Q�� 5aR�%t@3�sr��8Q@����`��vy��㉁ϵ.�
�GA�Ԕ�s��%V�]?O�9�U[ٝ��2e=�>g�ʱd��8h ES {]:2�Hmo0d7cI�+N����ey�º����ėHȽэ7~qC���b���D�!Tޗ B o���_����F�EY]�_|F�{��t�MU���g���wT��BR���зz���.E��L~Ѩ��]��lO&�A	qX�� S�0	��h.=w7s���6W��@3IDP����(���M"S.��W.���OO2��B���0Ď�[�r���h��'�7��m��T|KB5Z&�THI�����cR+,��j��)�����Ն>�ؒ�y@���щ���V�.%�aIF͓ ���ϽY?�I�ov��3���m�e��-���� �T{yH��y �X��%Y�)c	O�=8�
me�x���d]�|�)�;&?�&�1_�=��O�	b���}q$���B�*Rt��SΆ�U����ǩN��,�WuYR�j�Ʃ��j�i!
(yY�k)� �^��b�W��w�ÂvG�mk}�]��C��AS���w��U�&PZ�kt���7`���}^����p�i�� %���uz���� na�T�C�Hᅗe���FRoMS~�*l
�	�	т�Z~HyC=|�-��;%����9�t
�I3F�M��@�Z��P5X��Og����R͚�&�{���k��#�!6,f���vz���)of��9�P�����8=������e�Ϻ�.^�q<��߀F#olڭ
L��|? R/�x]�@��<(�͌�}2��i7�r>dP����Xǽ�+��8E���L�c��	�d��Zᡧ��B�H�Py52<�"�p���d����VW�B(R�Qگ{��/���X��P�jkK������JG�-Dݍ%9Ǹ�5��l@�;eԫ6������Q�l +���Dr��N^D�sK���±��KΝ��9D�ܥĖV�=o��wn�����V7�{���v��p��4��8"�.O�����Zt(48�g��e�2� 28�B�7v�Xn�;�^zӔA|&9��i�L�$�)�m҉�JFa�::����-*pA��t�H�~�#�6�P��e��N�B������Y�2ړ_Ĕ��& 򊤧w��g�?N�zn6�)�L��{S:�����?+�)���&u�ξ_X�5w3>����3�-%��;����@�WP\0�x�ڰI�9�;�n�:�\��F ����� %
�� � �_<_���n���S#�h�!|!d�r4��/uO�_�<U��"H'���'x�K���f�{���|�������@c�}�&�*p�R�!ڪ�:JHb�@j6�#��!a�(a�ћ{��DP���BQj��LC���l��Hj �3�`��{���ٖ������!1+t$�֣~�n'{k��n�v4��E\:�6l��'��;e��������K�����o|�ǭ�m�7�D�F�q�E2�O,���+}�����U�z�|;�����@T���D#����W��nZ�(B�UӕV_[w��qXہzp�a��K<>�4��4��B��|�W6cm}nD5��n) ���u��a�@,��lH�/� �\��E�ks.�T���Z��l�I��m{���N���4b�QЃ�(O~�ΔB�{�V:��{�H&����:��3������rsq�Т0���tロ���偠���@
�S���-+jO���T;��4�ń���]��$ ��*�f�®�O�f��"���Z��o
*�܂K?�!�Y��&7]�CZ���F�d��	;:�I|��!2B�a����-(7J����8q"�׫�eMGe�enخN��UJ�q��
�x��X�Qq$�h��N4���t_4xv���K�����L��ZBds(��@ڌ�l�F
�8�b��UGr\�C.�p����:8���g$>q����lE;��sB-�G;/N�x��d�F���Շ��� ڧ����.Se��!J�!?�d��KnΊvq�i��
K�LV��\o�M��I�P>���MV�z����)�)V��)u�Ä�VW���%	�����U@�κ4%[&C,W-��J�s�(��E�E�O�˭����w���K�ݦ��CX��}�@@n�7�Tn�4�"��d�^z�e'��������b��+ߝk選��G!X���y��S��J�iWy)$M�P]%�֘~�H�D�:Ѐup�+DEJ+=�ot����Z��pH�)�eF6D	��:�%�
l����n�m�^�}� g�C��剚�ؼ���PD��:�u`��4)h�[ �e�y�:�G]9E+#�8�o��f#(�|����Dk�Wԋ�ɭn�����P���[��._?�/��_#�s��}�p����'Q�S$�e\�K�t�t�RaAne�|a���RmyX4c�"�lP�=nO���Z#�Gp)y>����ں��?t:�����:�Ug�7Hl���{Ї��靶.nE�By�Qa�=�h�0�����.�1L8\b�]���y$z8�Ѐ8��Z�]���N1�7����2.�+t�+�~S& ��]��~Hל���EM�e�,퍤nv�`�d����� �s�#(����!��)����Q�7�?=�W�5����Է"�C�ɤ<�0�ȟPtȺp��)��j#�����I21Q�Ҭy����q�No�Q��;���(����"�zP��xj0�� ӣ����YX�s�Rd�6S9��(9*��͇��	aV��b���`ܝ��"Z6
�����J
�C�^tk� 3bᮑ�w������Jڅs�F�]�d���}�	��v�(0�0��d{��t������RU�]���� )b
]��-��i�I�D��&/s��Z��^���J�a�.E)�mY������J���*�ͻ�ʨ�v(E
�$	Y"��r�KB����߃�$� ��9i���՜Ɛ� ['#��.<k���r�p�ݑ�;*��������H�����~^x������*��iKC��RF��r���:#*wzLQ�!*��=;ˠ�쀤9���'Sh�eg~�����4V�hh�a!(��[��ZM@G�ԏ ����낦�v�q/��:zH�yKZX]�����G&���q��kl82�v����2u�[=(#Glob�>#o�$����"yPv�\ �`�����TUk����N��P���4}��u�q�U2�UW
k�lW}1��k&�r:{E��
�4?�G����H����#p���Zd=Z�ߜ^��Sw9΄3W�\��¬���};�J�Ju�k�Ќ&�f$���,��� N�1<��J�Hr�CmYa�fY�.�<U	��K@{`DC>F�g<Ĵ�lD�^4��"uh����_H��eQ{�����"&�Z��v�)��#_1.ͣ�1��U>�đҲ��u�Z��>�����8�=M�b���� �u�f5� �6��������N9�p�{g=�0�F���G2܂�$ ����2p�*���/p}W�14]S�'o.�?d��`�T\R���ޥvv���+:�_�un3R\J�o�����6��1I����j:�S�+�v�	����o@m湇i�@k=�o]��ښ�%b߷K�m����f���Scq<�������4N(��Q��A��q?,��ˌ����5�܋uW{��՗_�,}�^��S���)����/����upn̴R�Z���p~R����2��-m�v���Z���0���8V���0Ύ���+�qj�* �(�yU<����oR5:�~*�j���V��)��/�3K�+dK��O�L��`�NA����µj�L�Z0v�E����/"n���i|�VA� �M�I9�3r�QO��=��Fge�vw���^K�(~�>ECJ��4���ڙ�Q�����������G��D�^\�a)<�Q= �_��Rx�3'��H�s �e�\E��f�.��ʪό�QUv�u��24�,�$�iq��HY�+X剾��z��g��he�����z�2-�Wը�J8���&���Q��}��h;�0T�����ZOk�*'����(U[$��N�L�X8%��S9�%t6Z���g$j��U��^�lS�}�H�OxZ:ahr?�T۵N�G�.��Hܑ�����E�����4K!����iEަ[� s��)ؑ����i���0�����#s�?Y��{-�����zq0�-'B�NB���P	�`kõs�>��kWH���V�dSV[φ�Oڔ�'�U�b�h�/�@�aB�1K�|Q��u���:*���b��$���ԏ��O�'�ThLm�^4��Oؒ�ҞӜ��#Ly�9�����������ׂ�_ϝ�{M� �4���BT�>-�>q/lS�i�q��>���k۽�Eժ�7�"�i��/ h�M�!��.�唇MF	;�3����!�9'��,����ļ�}�+7m5o��S3��90
����W����	$�'> 	\Q�KI�{-FT��k>O \t��]tG��G�$����)T]�e������+2q��s%��h%Hl[A��F���� �i�T����vCN��'��|� ���xz�+9"҉�c��r�1��}Aj�s7����oY�o	�X���KW�RZ܄:P�!�I�"U�=jި�7;Imރ�t=t5k̴��a�X97�ӈѴ��p"���`�ۮ�������>vQks�K�CҲ+�a���^��EY!�甈�F�N���y8R�$�d��Ѕ]L����9��RV���	���~�#�~IR�IA��'�G���|��ƙ��,	#�Nh�J�*�����HO��35�Z�dUd�Xj��8��ğsV�b��ۺ;2�z��C��؊��m��G`���Ү�)M�'�U���!��&���N�W��GJ>2�fs͈�M�	ԌsƆ%ҝs\�����F2�/����5��:�]-e�B>o�~�Fܹ9�A����o�o�vN����7�Az���*lĭ�Jg��@����PŵBrȗ�x+߳�F�x.��ݪt���6�sCY�h�Q:��t��Xgz�;P�ym���֋�n�GN���Ј�Sь#)�r�3L�1���L�b�ύRg�O��DI��q�5=b�Vj	[UK��L0?&<�������+�`�X���#mڶ#�0�j;P�At&�����T6s�H�+�1s�@!�p�
]��"N���F��e՟z�{5��7�Ś&4��������nN���Yu���R���G������D��Oa����?9�{�v(�P���nC{F&�bf���k7Ā]��r�A�	j�Wh���u�Өr��Ղ�=+o��9�BY�(�u�>�Ogk��4Teh��Mj���[ߚ��܇p5 �[����
0��^���HeH�ߧ�����ټYf�z�G�\�W��+mx���eJ�Wq�x�P��l��w��1��s�2�a_��1nS��pyl��j����W<�G�����}�ę��c�G @�ٽ�)�夞��&ձx��y]�3A���� �~v'1d�s�q��\���h�|�K�Ih��۳]{��8]_C��o�p�~��Y���Ɋ.d��F�i�
�	/\�^B]}ޏ`\�ٸojR�0l�����MqA:Q��؆�y>��c+�J�2>�x���d�q-��cB%�~��w�K�:?�cy�t���L�,N�{䗰���d77� �+��Jʢ']�PH�=@lp[M����J����|���m����U��.	�Ҕ�!��FZ���J��]���j���[����5W��`C�ݦ�:k<A\�h	�Sԙ4犙A���4ip�F��q!e
r�O���9U�+��2ZR@P�E�V'�
��r|� )��I�۫p���|K��4�܅�����pB�F�KA �6mu<��gp���wuzyu�Gk�.��aV�^'������rY��:ĭBΞD/���v��-�A]Էl!��,+4��OAH����B,�h��?�{���(���9ʇf�p$������.³�AO�=�D\��YLn7y��L�e]p�ձ"|�	~�{���s��[D;j�^�,j�_�|ǡL����w֬�A� ������%�	����pK�e*ͪ�� �X�2�v[����SН�T�'rt*��O�W�c;�`�X��<�I~b~x���_9�<Iw��ǆ�hr+�%w��Sv�ψ^&��ůD#��T��գ{�zJ~��z�ME�Ĳȓ=?�*3�v������7�,�����g�0�ɑF6�O�Qxo�2�)bN�>�yƵ�,�v�IX�p��\ÈݗŽ�a��l���"��tZ��X��8I�Uz3�z���6h'!���@7�C� 7m��*$�E=���M{�e����&
�5�*��zw��?�bN�� ��(�Įά�`i�n%��Oj��|���+vC��:i76�	�F�}Y;�뜈��U^�b��B7y�E�Xp.!,e��0�*|�r���M��,���P�^c�8��$պ|��Ag��M�{P5������8�rF�m�+'+���6H崌: z��E=(%lXAN���q��_���1D����k���~��Ne��UPP�B�%��_P�!�>o����jG�!ag�di{3���b\¶�$(w��lD@ut�K��t�kA��\�U�3;��ҡw�ˡ�1D��	��t����l�J�6�Q����u���R2�~�b���g:Pw�yz^�i�����L��X��K�+��{�Cf�*�Ӄ"�y�����8�Ƒ]�R�V��B-�@}�'C#�Q@"��b��4� �[�o"��A�0�$�|���9F��%6���=�(V{WV2|���4��~b3�oB���uB��xp �7�Լ���չ�q�:f�u�6';-��b1�|��H>���Ѫڨ@�� �����?G�,��!�k��S���
]h&n��(�r��	�Y��ٻA�b}�H)6:}�4�O8Q7�i7=�Ъ��)�3?�R��Nʏ�	0c�zm�l�ǮC)�Z�[a���2�O�S�c�<�R������c�-d�����WϩK��^^@>^̡p9���_X� �_R����s}�Y������N�Q��P��g�Ꝋ�CW��� :� Zܖ�kqy���������b��ou@\7��hQ�k��D�:�=WZ	�bJĢ�0��!�?}m����~m�L5�-uy	����s��چ�78��5	����&A/DK'yυ�m��!*<���;p�9�����5��5%�y��� ࠃ��4�����*ɑ��Y��[��IW�������`�B�\aU|Fq�x1�4)�{�#�����<���V@-�@T6G��s�4�S�m�?�X�B��
ȍFyQl�K��$,;�����"�?��Z��ܜ�Sc�W�ILӂp�{�6�}����>H| �*s����4֜�߈���"G�7'����w�F>��3E���R}R:l��5�AW�;F�凱��҄�5�v�EkI,���Z@�ˏ/fm��2v�A����˻�j���%�H����h6d7�<���zI�s�ٯ��P���`��!�_��� ��@�&���cP�3�;2�Z��#ݾ!���?��+�w.�-��$��}� g~�)>~��bK-�������,����֡��R��	��-;�]w��k\y��K��s1���VͺR���~�cw��>�:�&.�
��jՊ���M�z.���wxo`�/nԙ\�2XS��f�"���[�7,1�~��΂����n���i`�l=&�[�O=.'��<K׼J�����e��'�, ��u&��	��c�M����ۃUN!
�o�Gnxb��@���h]�<o^e1��0��V.7K�"���&1�#�υi@���Z������26��Ѣ�3'彆���1n���ߙ�3_����W<�]�̸{��<4��u���T-�[�yC�ӊ]q&�s-IDO��
�#7�'���i�))�<ĺQ0�h��j?�bS�'~4I�L?��7�]qt#����VHl:��d�2hw�!��Q�n-�����<�<nZ�GԠ�!�M&Pb���Hg�}8>�g��ͮ��A_C����W��K�c)3��� �!���Wɼ���l�=��xEd3J�Q�gF2HE��9��h����L�/y#4��Ѻ`9����S�&Ą a�9rէ�r<<��e�Zv�]��z�7�P�Q��7�U�4��O����zw����׽d�����YMu�Av�����kL�	K`��)�D��>4���q��e��K���������@'�rh�?M�r٨�=���9�uY�B5j���u�Z������
SL��nC���1���EO��|e�^��u܅���&5�s�c��~�H��
8R&r�c�7�r}n�����
�����*?7"�E7�FB�XXs��4�j�J��Nr����E�/o�΅�o�'C�p��Ʒ��e����mǕ@Ɂe��TO���w�̚�yN����(��YP���h��v��iN�@7����Fm��xP�����@�'�w��GֶZz� %���v�!����|�su�8�^!U��WN�c �aX�}��������@��B�V��d�1:�~,?���g9<Z� `(f4L����-!a(镓tb�~V�p��b�\�$~�2�ȍ/�Xw�h3���w�w���s��ݓ����ټ�F*$�aB� ��i��2���KH��#7Thz��1g����w_�p�B�q6��A�}#�2�(��/WW�v���V&8�@iz���G��~���lk�ߧ��2�G��U�ʸ$��z�����fGMRn�gU�$Ht�0�ݭ*����}�Bn)ư�i�q4_k߮ A9"�C���er��@�-#��tj,���;��P�7phNٗ��oFD��@{���H%�V:%�*� �jrԍBsȉ�f�;R��j�YN_��a��}l:��i�ß�)�Rz] ����p��י�|���mA+�Ԛz�@Y�-`%r7+ц�.�}��,-ķjF7�ϡc�|œ�0x}20�p{|�oBh�wu���KG��-����1�
e�K4�p[�c���JU0/�̶���z�E:����[��\�߸L�z=�~�P����U�����C
�8�cGyݘ|�o�3�7x��fH{�� c������O�aa����TF�� r+�wLOQ��:�w�j�������D��w�d�a��a#���I���&��4�L�����F��d��n�MkE$R����`�CH����>z�>���2����
'��[�Cgc�@s��O(�c���Q�2>^b�~�j.�a"���fn�V��F�Cf�.���ZIþ�ep=�Q��4��?���9��n:^����(���6��[.�gG!��Kǈ�5%*
�އ�����f
Þ��@��tS���}1��fh$�)D��u�7f�D�*���`�'g��B�ri���L@d���ΎѳC��U�=6��ƪ����p�S��^�p�(a�gu�}o���_�S)NOgYaj���3"�J���,ɸE�H0k=����YS��mxq�EX�Īcs����eDv'J��oV�xBڭ�xd�����\I�F͋&o���W�f�m3�P[�������x)qPL�鷒��+�茿wH&l���y�:��C��&�4��`,ꟀU f���sG>C��t�=>7F�?���41Q햜K�P +W���:�O��:��������[����FɳU�>e��9�������>�&�6��^9C}P�֧ά�U$u�/ߙ ��&y�t��ӥh�	Y�3�ɠ���{c,���xzb���2Ց�伌���7���q��tw�q��%�A�&.�?ī��I5&E:�6ߨ����|j���v9�3�T�H��K�P�q%=�%�x����蝁\�����/�\��ô!Y�%�h������c����I��^��^�������䨲�j�K"�w��s��� ��3�$s���*F��t�:�1&�p�"6���� a9l�ރ|{�K�������>�Ӡ����q����0�A�+ps��澲(L��oV1��`:f�w�2��}��"������TZ�g��f�'��i�q5m4:��6O�����V@�;�N՞wb�%Љ�"�PZ����/0'1����S8�ǌ�f}>ĲD,��jd?�����X%ր8�.��qO���@��m��_��v�V��A~oF�^�vTtG&�@\�L�Q���>>&A$��{�Y�Ȟ6x3�8/�n_�f��Vz�H�]H��\�d�e��mƥ O@��C���h�]�	�[��|�;9�9�D���N��2A�x?)tf mQ��`fZJ����dE���Syͦ
�C�S�MO� <@g���8\�LG�z��L� �_i�LA[�%�A�2>�%\ԕw8�3|�)!���0�.NV�:����v��ʙ�(�����ה{����8iM��U�5"�p7�����^��RǒQAv�2?�iZkq��E�L���!M�~�i�l��ݰ6�ҥ�|S���AGRN'Ϟp�(;���5GzH6<��f �r��z��"���R.��=��O�}�m���g�(����I�ی�I�eWN�c�۝�҆n����*��v?�gpT8w>fsN�l|�d���	?R����V^a��"�gp/4�����5-��|�n	YK�K�|�Qn�o6�KM���h+�J>z���CZ~F[2��QBq�>�# �9T���.8mfW�m\�
��>�º��B�_<�b�>�"}�:�i	|E+��TlJc���(����K�l�X�xm7�a��,�4fz���0�UUi�
>���Ȟ�g��|�C�ec�с�馉֊���Nw�M� dͭ.�t��u�^���p	��Fp�]����Յ��.��p?Ӻ�$$#"���B����wD=e �Ef*Y���f�G���Gx���zsR�!��]��ñ,|۩֡��O���"�T%��ZC�=�s`D�e�ic�n�2�������^�}W���^�wu�_��+ly�fE0c�B#D�o�����d}!�����c��j�����w���n��qi�Ή8k�S���twMƯ�C�9�0��_!+!ί��U�Z���lV�D�]�d
c����1�h
�ǀ���u-flq����9��'�f�q�D�yEp؍T��_ܗ�^}Y����!�)a6$�S�1N2��fӭ�uI(��f��Y�WxȯvX�%}p�����p�-���O��Ԃ:�C����NU�Ƕ�\�nZ�/Khd�8s�.�`���N�~�@ գTm3��n��^EM$��H�?���o�vl�.|�	�,Z��t2Tk�_�N��\�"�֔䆎"��S���lJ��!��&����D�z��2�k��2R�(%�Ǌ��@�{���>�x�l�� ��c��nN���2�/��mL��*��E��dj~�V��I���:|2e�s�ލ/q7&�n�P�0G�2d����Ҥh����
g�Y����Zߛ��U���R�t����<$uqO����5xߏpI]�DT���E��q���MŢ�������[�7t�j� �=���#��}��~,O�|�b웆�����G���7֣�#�7���sFW-i���C�����1R)���s�&�]��JRfd���&tQ"��u 7�A�-KV��&:� 	��ʣ�e�Q��È�ʸp����5��k�/�:rN���,�l������� �˚h��0Z���1��5����/0�A�uP��g���۽m����r�Ð-45�5�W}`f��m��^���q%��� �Gı�r���.3��y��Uu�M�c�A�ǀ��h�!�2y�M{g��4�Ar9���D���/��9�S[���q2+���.?Ç$�Q�t=�S�&�ʜ��f�﵂��;�d<�^h?�	��s*r����ل"}J�����o"���Hu���Qڞw�󮒴�*8� ���Z�&���
��a�tFh�7��X�;��_V���y�����Ɛ�n�7�}W�,�c(��9,!�q��V�ASf!�=��N���X�,z��.�r����0rS�Y�+%]I�.�k��2��6NH�GK�U����J��]�����A��Y00��sZ�3�I�~?L�7�`�����ʧ���s6��
��t"S�A[�&���I>�~��_"��Wt��f��� ,#u�����S�
-�n��!]�����¬q����VDa�4Hn����-���̲���aS���Ǯ٫�������j@��k'D*����FZs)�0GiWFJ��̆�Xs�,��L�k������XJ�h@������B�b����^��7��U�
��Qn����{�\n�-x�EaGw"�$o����x_��"_,�����NؓdA���=Ć�7� �w`��(���-,y�93�d����Y�	�ft(Of��D���"���`aN$��m�u���o�W.�l���Ⱦ֍h��ڤ0�����j+�4�8�#8n"Aޡ]x�įӕ��zOy��_�`��[� ��͠��(+jQ�!�'_�;Y�Ow���x:������عM�R���U�U��"�\H7�ȕT~M樂2���|D���cݺz�&����Z�����f���a{3������� ~���kl��_�	�-7�vq{�
C7�bC���=u�N�A��H��J�Q;_ǝ�d��V��4`K�èwpǧ?���IcՐ�� ��6}��m>2�!���l���n�f�1(�.�Hf
/��Z7ū��@E�BInߧ$�?� +f�zn�d��&vs'�;FH���G���W�\���=.K���7��i����-��K69���������P���%����W�R�/����Ᏺ�l���	Oj��|ڼ|�|���ȒC�B��7��-,�U7�K^���_V����ȟ�S��ѿbay'��vz������������C+��b<k�����¥�H�9t�h]�����Лn�I|e�O�(G !N}=�XN�j�(y;ͭ7u�?��_զ>�ɗ!�^���Z������@Ν\2�����|��*Uӧ6 R�-���9V��^�rW�dy���O��2\������RX�9�\�0[M�@l���49��l�_�V�����4c&��	��Q4��9�VIě��*d�ڟXʭ�ϲ���
mK �q�y����pε1���\�U Ӓt�_s[�֕O�C��pn��:~�&�>I,/��З�����7�#�jL�ҡX��N���,e�%�|m��V��;�
�Ioq�-���ST~�1�mϸF���^q�Z�0"�2����֏@o�{��.J�T�x�szc�'�����%к���ZRc������!X�B�y_��� ��t�yJ�6����#{��6T�my�#odާ���G4�I�̺V��Pa���(7��|���bC�B�v.�>}�Zn�!L�/mHn�r��d�2�:��K��#��z�Y���!s3i�"�/e��vU?�����D}���J�O4�����6���u�f9����z�Yc9���[L��Iz\h{�?�1���v!a��eU�,�_+��@�X;<�iA��0K�x�Q�0<}�W��{�i&KFKx),eR���r��3s`R$w�����e���|�%X���1�")Xd�v��P�݈����Y�l��K�/)4V�)���R9�K��g:��4��]D3�I�m��Bz���OD�s��i���5/VE)��'�")�%ᔍg~g*�� ��J���x��3_1�#Źf�rB�SѵZFÇ�����&њ�Yv�k��+n�]���#d�ښ%nT?�����"������3�vvi����B�
��f��I�q)�p�����Z�W�3���,+g�=%����PO��>�D�W��mK��K,Ϲm��QcGc�@1�Q8#ELo�r����g����6M]< 
6�C���`��WCj�����m-���;צC��|2���1* w����AW����Wʯxho؎��������ɖ�l8�'>���HG�и�]�m����^���F(k]}_���lg?�_�ރi\@8)��A�̒ĥ���ů�26�U����ޜ��KeEN<�N��хl�G�/E<�N򫃒����޺p`��8�"4j����*����8�T]!���f\�'�ş��M����I��*�մ�N�a[�i:�ap�в0n�[i�M@˾�����@���s��V���Da����\�|�&S��B4���}��*����T��c����PXM��6�p�$�õHD01𣲟�:l��NF�d$�St��s��>����Jd+C3�{w��o�`�F�6�ƥ��l�%ߐ�2�ն*���� ;
̣6�hN�7t{S}�YL�tK��5��P/:=5��T��Jژ^2��[=ދGzX�w��>����"]���u,���2����D#�� w��qoq�)V����2�_�	9죽LM��pؽB��D�2|#]�\���B+�sl�Tܬ/�Ė���Rq���H�'>�!z<�B��}�+�Ŷ_��EV���э�kE}9utc�0���
��(�P95��9n~
/_2�}0�!Nx�� 8)�&�1�_uw��o��W��Jl2�� �q�O��vi��,ॕ��K���k�D�ہ���=zy5��	��r�*ӊ*A؍����1��ȝ*4Y�D�������w�������e��`�
�=��;��]m\�*n{_v_��\$�T�K;����~�OK�.�4@C��6g�*~���3�G7��c�PU��6JhJ���:%��^v2���]W'.�YR���xV"iYa���w���k�ð���(ݻ��,
���+4��2c�N������,�iDs�:���6)�dIn���Q�@�l�]51Z&�/��>��.��$�Q�W�"r6�@��EPs�x)�<��,B.�0��OZ�h֜�U��'�o7��M���3͵���R@7�b�aӠ �%�6�$WwK̵A�^��arP�3l]�D��>ك��%7S&1S��M7�f�(Z@�lv���[gK��E�C�-���)�QS8(tcD�@�c�"��d���Ф��nj��X�ǳ�Qp��=�O���\7I6�k��w�.��2�����I�A]�%��Hl��j�8a��ǿ������L�\�l�Ӂu�Xo,�X/y9�=h�E�����v�_�Ў�DU$SQw�61��ȴ)��{��=�<E%�P*�y�T������4Ssj�.KοAV����a�<��@�k}&�!+P#�(�?�E��'<߷�ا��u�Q
%/���'.�������ݯ����!K%�-�1�4��h6VY(�Hb���k��p������aIt�Fl�l�������X��Ih�%_��Z�?�څн�W��_�K����#�{�y�Q�5��w������&؍`���H���H�HXw�	��ǝ����Z���#؆��Ȟ�k."�ٸF��e ��(��D��)Q�*�sԯ�Sf�P/�8������|5��p����,�^�j�9� �;�a>�K&H�^g����?�n�ж���V���\Lw 4��ʤT�m'��P��m77Z� ���f?� =��0�k��@�@8���E����(57��u���ATp�Ne�e���A�]�h�d�θ��7L=ޔV���3xr<HK=[e��)��P F�Î�%�Ҳ���r�F����!�s�\�!�+[�C�Fi���MW�ċ��Ҁ �K��/�:6�ݧj#lh1@��]?>���E���?�'�E�:nK�l[I���䈣��֣Q�����u� �fx<%�b-H�j��W<9�<@�U�}]\?Z��&�a:��fǇ��h�o0���wQ����sf�ŷ�T�t������t���Z��cb�"���%���2���]SE$�̏(O���wT��w��Oڻ���K�q�58�-���g�&����`�����@E����*��(���n��/�#TP;�	AJ�K�"�0'�ŝ)����G>��f�����7��A�>�����t����gBad�	�2BԪl�r��U~Z5���
v��	��qZ$	�3��Xq��׹�Ҵ[�ws7�����.1f�!gp/|Pk�~+W����J�kݿ>=�F^��y\mq�~��)�����B�Q�\ZA菂�MN<��HF��^��<�Y	g򘧉9���O�Cښ�2�'��*�[4}p���A���pM�m��B���d!�ع~"����hګ&�`ASV&T}�0h�ߧ����)��%��G&<����]S�Y�3I,���n�5)�����&��g��Z�4�:&S��r�����a�& �� �Q3]^qⲗo֭��੡��0<�����7=�ˮ�r��?����?[�ހ��C�B�#�p����Q9[�Z=�aL�7�$q�߾����Z�D��ݽ�|�)X��G>_��}wn���4�FL��fջ%�|� �bf��!R�6s=�*���9W@J!C0�PPS(g��w�o��k�Y��@W FoU1`4�� �i�#~N޹�mOE:�b��B��×~�H�e��gB��,,o�y'��7K`��h�����P���"kXY0��"�������CD��-��������%ԼUjŲJK��!��\�UghmL�P�;}f��C䫨zDt�ёDa�+�;��x0�b)^2���"�zl'�_ኤcp q�&�AS���N�`Cc��I�u~���3�4����?��!&���D�V�����BJ�F���))ގ_��|�<b�����x��ځ��5���=�Ba/������v��]�`�V^�\a��6�Rт���Z3t��_8?��F�x۶�|�ׇJ�a^��GM+N�,1�FF��읛XD�9�7HPXU���c4�4��KWM�y���[�ŤN�����	o��-�f�u���bP:��zQ���&�~KU��&C�S�a�Be��.��4����E�<��`���n<�� P��N���[It�)�jA�~~8vjE oA^Z���Ӳ����2����0��: dwr~�i�GtQ�Oj�i_��$�I����_$C�p�9���0�;^����<ѥ��r����S�0��U�C�ő+Ӗ�E `B�ɣ@~��� є�[�f�@O[�RB��������rVM�VUMV�d������M|�@���R�{H�c����Y=@�sC�|���d�.sΎ8���i�Ǥ�d#���Z�9>O��E��|\x*[�}զ4����;r@E߲�R�()�5Zm���n�y��ɫ���N���G�j\�c�}:���
�e+�;C닊G���ܟ�֭;�/����׉{(��aǡ���XL����-^C�$�HZ���;g�`9�n���פi��� ��o+T4i�'��k� ���*�k��s<x;�~5�R�����/��8z���|/���@pe�&�*S��{�J���2��$�q���XJ��¸������P�6ɇ����@���>agFI��x��� Id�h+C~g���?�y��pv���8S~'�NK�۠Q?4M�p��&�#,E�����-@�l�Oׅ@�f��D�cd����K�|�G���J���炂�H�iA���k�^0�FW�d�IIe�����۝}��	�bJξ�+��O�C� �`h�&��8=2�����b*����O�+Ԧ��S��kI>�����iH�M�>t/����+0Cr��k��zN�ϾZw�#V���cR�h��;C�l_����zi:>�N�kyjg����!����m�sT)��q�������Њh �i@%��-�����5^
�bSŻIo���VQ��Yx�̷ƥ���-�Lc��Oa'��5|$�
��'�?�v��E7��O��b��^ެ�þS�΢M�f��g�@��?n��b��+T��)yDq�a��S��D��딁�8E���Y�_��` A�Uj�o��0UJg�!�^Ai�����U��c�9����bY�w$-9V��jԅ�Q���n��88�@��8��O��Ѓ��>����4���s���C�q���C�ʽ�6e6��]�o�����1��Լ��s���^j��ȶ*|�ّ�{��`�\Jf��3ש�~�?�Ȣ5�Z���~����Yh����.��]O-nMK�rA�O8��T_���.ҍ:��R��֖{1��q���p�Lm	�@�Y�ۜ�~6��y��!�{By�@��.c�xnw�<������&�3�����ׇ8˕��T�R>X�zyP�����jFE_�z?��� y����q|IY�[�!١�����;�
E�KL��ʽ�d�0��p����Q��TnMϏ�mљ(����
Eȍkȃ��s,�]���C���=�G�Qv�$����G�T֝k�q�1a]`�V�w9�6S���h\]�_���z��/r]���-C�,x�Iv� ���+�S�� ���
شٮK}˭�p���$K�[��BA�d�fVk�EaBs����	�������^���4Y�{��֜�y���-3�4��/�x3/G��H�k���~�9i���&%l0hԥ�4WbgPs\��϶�Q����d�!�uPaE4���Tg?Iq�/LR���)�.��D �Ыd�)�f�$ssO@K����c�`y�62�m��!~� ǧ��ݙ��z��s��<�l$L�ެ���<St�m���Td�����DܬǾ�O6><)����y���1)�L�㎕ø���?⋻�zw�Tϋ�eb̈́�^�����L�F=EF�}�A&gt��<�)��~����v�$Q��r���L���@�:,�n����k,�k)�(HB�Ŏ$bpL��L�^�%��.G`���P���yT9f�1��l-�M��Q�;��۵���D�HIVA�VO_�Ɖf�7U��'z���S:ͬ�,�^.v��k\a��waSW���#U\�Pև"(m����m��	��R�����c�=�9L����m8��yӹ��B�)��<��ɨ<0������=��y�����N'?��q�l����]hPS ���1oq�l�*�vXDh��7�������~cl�MAV�-
��1)���MO쥺�w�6��	p�v�9�y��W˳���*�[�.[M��ϡ��n��KqxE�X���DJ� �������A�<�\����E����z�-�o�m��W� �)����Ls�%��x���G���ҁnq���lyc�;��4�*ܡ�Zk��W�o�ޚ�F��˵&1l�ߔgms�=�+�~�f�ÌY���|TD1~ǍGG�'Z/�e���KZx��qr�U1�һ��y!�ϰ�U�&�R^��i��4�qfD"=�����z���� ƾX-v?�D8�j�c�b��O��%:��/|w"v6	a@�6�s��	�xD��?�v��x�~� QiS�=kq>nW7�]� �?��؅���O��t�"��v�H�k�H�.�1KC{@"��[�\�� �6���f}�u���_'8-K�&��4���߷ˮbO��������wpȾAG�
P����>����]��+��J�P�+��	،��n,˰��`��<2>7�Sj�jbG��:8U_�@���Ǖ�qF--���G�ic���;L"(�<t7�e��3��%F�6�Q}p���e� X����~�7*�γ�H�4P���arl�V˫�旅�-D����Ek~
ȭ�h�0ld�uR����p�ϩ�T,��f& �ۚ-��[�HYr8I��҂��,����]�Z�8>��O��XN�6K%������iay{��33�~����R�$E���>9�|.�;FϤ�>W�C-%�}W&����q�5L8�{�c��3��كu�!n'�!�g�­��˪!�@�t ?�y3Q�6+���L=��6 ��4���L��K��)}�����!�1d���.�j���E�o���W�����r�k'G��l���?P�2�p�}�W��}�d�9S��7)=}RB� h�zn��Ak�|�*b��7i��s�X��.F�������ޚ�Z4�e�\쉚�H�*�<d|�;7����Y	�<��Q]�DD�DM�Ո�}���?�23ܒ<�3�_Ke�ù��f]�'م4sU띬I�C��|���b�D��|�D�3?x�=�%��4���î��v�����X��7G�;�r��3����M���]#+���a�h��`x��У�6p��ox�#�7���X�������2�9��zx�B����6���ع?���/�;��=2  m *nM���.]J2��Nz�Ӹ쨆�O�=��;���d>��-���
���8��$������)�	�[=�8��TG�y�����+�욾#�@r���k����^��F��M]��~�&�Zb y���׈�|���}����ì��ԕ����x>������po�Ag.��U4"���I����'���h1t����,�i��ny�暃�P��NM�};�EOG���	fzՑ;��M�95�&��/3����iu�
 O8��p �V��Nf�d���e��XJ�}gRg��mHo���B�B�؂
��]1��ck�'O=d�~��~#�j	8TR��q�,+����r��oN�$�F������ \�&ŧ�'uW�7�3+�6����P����cX8��h�B���vǂ��3�*��kA�-?Q�z��t�� e���r��
j���ɸ��Ii�V��܂�!�֤s7���_���#~�J�'���� � ��L�ӖD�qK����/A��w�`v.!,�|$���9|��uDx�l�������!�8�=In�z��n��ׁ�7��E]���8
���W�Ə�y�yCe'P�]6�����wX0���"�
�@,��R��:|��g��ҳ���|nl><�AE2N�y��.��O�����Wo~lM����:hc%śa�q����{�֌�gx�����Y,��?�N�[h�v|��r��LL7�Ư`�=:��Qٟt��ô�+7������p��B4}��#�p>B�پ���6AUNW���O4'	K��ɔ���`t(��V1�@E���X��?&�qQ����o�����ʚ?�Jo�y��l�C$Mf���j���M�:^��hId��n��o�AՄB��^\f�*���iP�4�% ���#�OV�� �HmLE�)����������(
 AoTv�[��F���⠨�h�
�9��j��'pڡ�{�)��J���P�x�A��f��h}!��|���p8��d��R��*Ǧ��F�n��l��_�=�����Eѿ�i�3�����XZ#qj�{ߴ����q�����!�8%���Z�t��z2�A6QC7h�m�1�~R(���3�%v����T��5�����N3Q{Թ�q�T6O��wLҪh���5�[v `9ʝ�j�bǿ��fx�	o�]5�I�&׆����ٔN�ю����웗��9w�.�-ˏ��MӄW-��:P2a�$����y�<���eh����?�8�m�o�*�%?͖?�b�8�S��:��WWG�R�%�rK�6.4��o��L;���u�ù�!��Va�ֻ㠗�{FB�^�ǣ����x�3�_�^9=gN]�:^�/��st�Eyx<����Ϣs2�P`Q�u�(&x"���"ύ�;� �x��I��F�e���(P��w��D��U��s�
M�n�Ln7D�0�:/��&lD���ON��i[�Pg7EfC��*�Qcj���h�b�l�S���}���ed�ڃ�D�rA�:<l}:���#���$�S��-g]}R���9
�T�q1z���x��������ƺ�i�0fm	����H젫x^��<�꾌rO�'��ѝF�����X�8�d8��E�:C5�^wp/e�9�]����kwvm�Xq�ō��0}��m+b��N�"8���g�}���dK����&� ��CR�#��]+�9�V��2F�"���k�~M�'��n�=�]�;�,w�ٽ[F[�Dnzkʓe��ͅ�5̹�_��U�c�1(A~T]S������mq:���e�ֶ"���+ó���l��Gw�r����>��sTp���.P���k���%���K+%�d����O6󤭪�Q�l�/&\��T�-\}��g��0�C�,*(l���� �@SFKZ���~ߦ��P�SȪ`(_�׻�Q|�n6�*r�-��#�cB�n0b�N�WR�$��͹m2���+��L��/(�Ib�q���(�_�I?f��s)�ٶ���?_�MVʏcb�?i}`IU�&�۵<[&vN��n�Df�,;�n�	Wg"��YcC�Em�ɋp�Gt�oh���hL�`З�t��uX�XI������z |�@#��#�bY)�i�pD��� #�k�_o�D�I7c
�\u�V�������w'+2L���ݐ�̗n�:�Ix���`�'nl�1�n���`9l:�!�&�G�L���Y��<j/�b<�~j(��u1)��~S^9�Py즷�f��	�,���A�_C�����ْ) k-���E�^��VoQ�T������N�0PUvּ�z������k}�*i��_�ea��u�p�x�0�o�X�|P]�q�;��S)�$�r-��/��@�$e�8�-��u�R�l+�'?��˨�e�bS.���&�iKq�F=��͂��9|�h����圳E�uau7z/ˠ�3����/�F�T�d^�X�!	����"X�4x�������#0'D��#Pu`�f"VO?�L�|`wj
D=İ���u�'�/^�_�}�<���� �2��j���Z|}��������|���@z��eM}�m{M�#�½A�ݢey*Fq�D�E#�WJix���sN��ÐM��Ǫ�(��y=�$�)�픆�=���z����.�k��a��'���deA"�k���Ng�GW��juY��2���ΆT�67������P��)(�>�j+���)qM�K��G��.�"\�2�I�P`�AEv�)4�<V(ڸ�Q���~KtRi5JNh�fS��q��&'����\�!�唻_w�����"2�\j�z "P
t�?�I�����ؾ,�A~W�	�:�lY����<]���}|Kv�" x}����3ʮ�u��{gyh�<�x	ivT��Z���L��������6���]��?
�~>��ߡ��(�hBH���s+���B�U.)r�oXn�Tbs������נ}��e�1���C6�
G���E�H�����xP���e�;�r��X�0��<��ܚxƼ���9��	b��tRA}O*(j��7��v��P*�y)C.��gݗs����h�^"���x�P�U��x�S�	 �7k�=��}3����Z�8 �D$���(O�3���jϹڕ�J��2x��J�m��b����ߙ�BS��{/��፠��H{�u������;�f��&����q��EY���1��H���)�9%��I����f�n;�����a�<e�6^p�e~�8p,��}��UY寧<�p$�]d�+&y�'G��ip ځ�g�v���K�)���(#GF:H`2,&����&�M�4��f�*��s�)l��L~�`F���,b��Dz�m¡'w�~'�2n�/E�i0Qc+��� �>�1�Í�됹jt�Qi���U:�4���D�sTx��s|�I�C�a�'�~/�D-�_�R��X���d.��4?�'���I`�����%�ķᭀ�PQ۷j�uOiS�=^�1�ȗ׻+-�үU}����0�������t�}���:�j�"�gx�S�e-< L?�םx��g����lyѥ;�dz{����Kq�]�].)8�C�������
�p�����k9L��'���4�	��҅���x� hP�0���+�i�ƩQF� �;��q9��M�H����	v!5h)\��h7��� ������ϧS�gp�!X�D�YǛI��㢯�*�'�V#{П��uz���zV!�����C��jZq�P�������l�����wo��S�j �����ux�V*�{=my�`2�wzC*��72�xwړ����UޢW�,���e��3��6���B��]��l#;o6RI,����%� ���M!�w{^λ1��I�����4mx?R�^V�w�"bϓ�\�P��7bP^�ߤ�Q���m��4ǧ�*z.�P�nvQ|����㚫6FNI�QT��?4�q<���	O��2g �X�w�A�N�*��;��j1�Ǧ�mt�����|Qr#;����X�_V��ŋ����s��z��U@�Q�o�j0y�a~���O��<� t1'�Ħk�\������eP�s������X^�

�Ɔ�'����\(t�k&�q�<Q��m���5%o�ѓ��(k�����2�A߳$s�~k���1h��=E�+3��o���g�S��T�~��4kp�4�.��d�� MGU�q�T�PX���Ô�7p��wǖR�2�u�;�`��*h8�&/ࣀ�e�V��:
ʅL�~q�l|�aq��.}�c-]1 �9�4uwx�SFQ�>~|�
���2�U9�Z��$��ܵû�PE�3�V+pj����]����� :�[z�]��{�cI��=b�C�9�)�%��k�c^�Y.�B@~`%��[�7J�{"��SY�P��<YD�������mQ3*����<�`���L�i�k +m�)v��|����%j�2���:�aM���F��%��f���|.	$B�݊��Ǖ"�,���`U�	h?``���-���0c�z |�8Zty���W�Xli�"�_܏�k����d�{l�՘�>�=��H�N�5G�� ���]se�E��O��&�Kޏ�������Hb�41'�%:�B����?�%�Օ���/U,��u>��^(�ɬ$�EY-�w9J,�y
� �Ǟ��>�o���� �:�<�x����N�%�CN�iJ��y��_بp ؓrx[���@�GB�5&�S��Û�N� ��M��W >���IC?�O@Ң���t�fJ����A%m��CX��v!&��j�:.ŀ_�Ƙe&��LQ��k���n�Ou�#,�q�[���AxeCڸ�;��H��a`+�C���e6 K8@��by��6�|��Njxn�R�F��Ѿ(��A
:�|<��x��UI�_yC��釔O�P�S2dw�xe߻9����ez��,/�(��T�!�N���3�u�ʌ��QX��D|ڱ�.Kui#�,-��� tȁ��D1I�/��H�F��	��}}\�����O2]��yR�p0 ��^r[o��g'��rh��ƙ���ҽ����uqO���m�y͛Y9�6%�[@����Geļ��V+t���j�p�J1� ���5���&������X�]f��s1�aJL42��D�i�r3��<X&T������&����Lh�w��`����f(�]
�fG� ����l=�:X�aW�M5\�e!���4�20s�[��� ��դ���O%�yl?��H\m����jZ	L=�mg�|�C�q������ʟ�����i$VjD�8��02L���U�9n�2�ހSX?���S݆31JF���2)3�4@�R�O6U�g� �A՛^�X�D7%Ff��ZZ�}T��_��T�ي��v>���4�Y��$�>�ۋŇ���axd}���-����d�{�b�50�q�ّ��A�9C,猍'�E�l��3ڂ�)X�VP%@�:�h��޷0��6�]��1K�/��l�=8���@
ϯ��~�eY��6]gW�M�����mƳ��#��a̿�Lr����&ghbI����m��������ϒ�8����[E��V�,�d�c��Pa;����I�֣����:��8Kq��e���i\������$�/�d7�A�riƻui���T�5��^���4m6� ��omj����Hit!'^{����V�c<8Xqk^s�Lm����ۭʏA0��iI��E�\~�5*���U?�33��>��,��:h�
*沭-:G����C5��V�I~jC����w���n��k(�ұqX�I�|��t�;]�]�%�g�(q��l1��|9ٹ�#�ݪ�j	!��h�o��v��&)�y�&AY�/���Nd����[^�;:C�S0wn�L�rmL���	d����o0���g��5z[C��w?��Q��X����%�e��{p�K[�0h)%��N�덦G�*-4c�=��-,k�`���[��a�<�����5����`́֊��e|����q:F��[Az�Q��lbOvU������AB��Pʥꔨ�i�G��|�x3�������߁�\�y$q���g��r�m�!� �f�0��9ɷYy&��n�vhR��|�CkW��������� 7�����w�U�����U��tQ3e�>�.?8�IU4J��o6�Q��T��Xk�b5��^1���IG��'7^�pO[��NI[��&sD#�(��S����^�Z
Iȵ���-������t��u�jtO� �����֝f�#�mM `�����Y��&�h�j�(ͨ����?�hl�>�Q�r�@.~"���8Ap)g��>���AW�����O��vר���J�!��� ��7���o����.9�Uv3��&��oa�+o�8p0�O�]�~�T:����z�����|,M �gB�6��6����F�<`�tm�C�m�a�v�n�I:}���kZh�����p�>��BtS��LM�`w��"!��by�����J�&�v'�RsPim��*>��yN �ly"�s �*@����e��ԣT�z��,��Ӂa����o���?�I�=űQ��Ɉϼ$���Z�]�hDY��/�A�pM�U^Y��=���a`�#��� �Bz�u�[3��̚%��=}o.�ڲ�	��=�._4N�7������!`�(��R��81��N'E�{�?:8������n�H'&Uj4?9�������O~����
DU��Z���責$�p�9a�������5�cf�٦q@��\ɣ�j��OE��/���4x]�Q{�C<�ӎڌ|+7�K��܉wR���.�rƒ��8���s�~^=s����E�8E�vM�3Q���$��$+�&Fe_6O�\Gah�!���"k�A0xH�n&7`�y�5W����W�O{K 8J�j�"�l�b��c:���E�`��qV�@���id�_�&�-�}S�����P�WA��[f�!�ʵ��<���j���$��|$5�,��� ���,�8Q>��/�v������
+ � ���[��0���t%N�{=�>HE��^��t��&�1��BY��v���6�$N�,�0w��|�L��\���O�Z�*��?8���{���v��1�g-�B0���LЂp�H8�^��9���N6�Z��E鼩��D�AH?İ��$|#U�������Ҕ��@�C�c�/aA���=�i�e�j.7'z��r�Y?i�R�1�b�tX��<��;�z���G���{8���8+�p���4���έ����<�L��b�&zO���+�o!`Eu�4��9�|$FE�`=3}�p�Y��C
�F2�!S��\�!7��,(k#�y�}a.�G:���!�Bq��v QF(���GP�`P����]��ۤ�+{בxOΕB	UОuu���zw�T��w���wÍX�؂�9	Dso��ҡn�R�3�����Xp��$d�\9������\&��J�^����JD�(���ូy鹈�[+�Ko7SUd��j��{��ɳK3�,�.��f�qǺOSӐ�t�Qȋ`lf[(x�S$�F�e2��*ؠY�${-�����Yۣܴ�u���#����/&�IzE�!���s�����օM���͏� -s������%�ՌRa���7��X�\���HX��̡�4��-oHǆ_^d �(A�*
��|�ä�3�k<9Y��'������6��3:G*�gbZ�x�M��mEQaMW��{j7��U����\Gs���2��enR9f1�N�/�����`W�X��x�5qv�kX��!&���_b��9�{���R�S("�ͯc��/��{CO>�y�7��=0
�t?	��چ�K�a�|;z�z\�\sM3�h�^8���d1_�{̅��Dƭ'��A�$��:�2����V�h�$!lLV�2�#��䖩>d3xZ^(ƻ�g������n8������d�"���a�兀�l.v"��B��X���T�R�X�&2	��}�Vc���7�M8�R��d3�&�c��{r�� ��c�Y]�v�Z �(���##&����eԓ�/�|�K�Kn��:������) FX�~!��Qo���V^lBQ@Xصm�n��~-�퍶�J�s�
Z���a�ʄ�X�%!lTQV2�>�+��IΰSt�f3آ��A�Jp�����R������AjA>�W#�&��D�$9�/~a��	�s�t=�Tmr5P�.�����6��Z�bM���v�|��#����~�K)��Փ_<r;�	+'�o��������ȉ���=�a��B��f{=&KtԻ�(#�O�R8:���I�h�'�\���D���Y�f} ���8���L�#\'����Vw�L���G9������w�iZ4R#�tB�����H�����E6���i,��>,�`��H�9�`bZ�tۅ\St�爂QDB	!A��t%¶���׏��C�6��}�ZbR��R^
P��<at=0Æ���2�ց�ή�)��6_V�O�^��E�nⓂ2�W(:�5�丬xu�X�{�%�C���\d	߫mC��<#�� �F3QDu�X�A1�+���X�H�E���*���&���;�� .	XF"���	�w�eg"�R�Hn;J\XȆy�Q�]�i	|�PmEQV�Έu�ݾ��\m1��%`�2����Ȳo�F��K�ɲ<pܚ ���X��W.���L��K���:���n�W߫��)(@�؎�A8\<�-`դ╟�e����*��Uq��x��#��3���T��' ���erz���ġC�3��p�x�_5�)\ Y�n]���u���+��!��a���ks�J��&ݓ�Qű����n"s���_׊3�DDJ�O���{�#��(���1�vu6��46�^�YX�En|ӵ���mY�.��ot�2|yU4�P|�Cv��N�4��t�m�9U!`����H��)��h% $pWE;��g,�g��\�eX��
��Hĝ��
6��`�*-�F�	��YzU�ʇ����@?B�X�BJ�ֽ���� �(�f��e��dI�(U4i�r�_p f��m�N��>�8(�d����
X��Z7*�3�Z�f�Ӗ(k!�'��n�?s��ɤ�0E�]3$xZAk��n��O���9H�b�J !rW�ف��ш�ӺKW��q\�X�*�\sﯶ]4.S���Uo��=�+��A@�:f������JA�!w�0c��N1��[���$PC��/�]�.��-W�/�^����Jɞ��R�l�j���ȏ�PQF �`�
��2��u�(c���!�u�I�Pw���G*IP.�ʯ�!EE��ws��VBZ�R��a@zF\%r�D)�$s6(8M���G�*Mc�$���V�Sxո1߉+qb�l��3P�����d��k��q�4%���&����\���ED�/*�no�ҹ��ű�c�8�j1� efR�YSL%�C�A�nI��TӢ��% �����is��?���Գ���޺M '!��s��Z.�.'yx#(�ټ ��K�f������n�y#(��׊���`"V���(�~�G���w5vW��I��'k��8���r��u2�1��!$���uf���m���q�m�E����}o���~���i<�%9]��(��a'G������JS����$�JSȡ8�2��g��O��CL����q�K��
�����`�r<s�%�"���p�D����T`ı���[��.��AV3S��Uߕ�R
Kz��V9 {���՛R!�|�^�>t��fx��Q�/���=@o�tv�w��� ;j8+� p><�S-0��x��[rN3��3������o˹ z�=�>F�m�אx��ӑw��"]�����^�W�~�(�c|M�������:V�xh9N{�gb��U�_����v��=h��fO|��1��l�1�S,�-�_��s���X�<㎓]�C6(�-Hm�-���c��W~��<�7�����s3�u��@x�;?�^.t/��L>�@(��b�U�j���/[��e�-�@nnA�eT��:�ހ0?{����JV���.�a)��߸�)l���/�S\�3
�!v��,)����T��{�|���+�轁z������'�>	R$���nK�ͫ���V�"b� �����iWr$~o�Sl}�^0���z�H]EWh���m$v�. �!踇Cl�ե��^����6�(]J7��8{��H�L��x�8)��`�|~j%u)Q
0��⡄ҢG�f��&�����M��P��s�W$�y$*:�tiw�sL0�/�E��팍u���s_~&bmt��h���8D����%��qf��b�	�kxjJ��(�-�:��R��H��g��ʯ��O8�x�}�D�+f;��.�rQ��O+�g8���>n��|a�W
�/*�g�М4�i~_d7��cҧ!Wv&w��,�<:�J��KQ��|�Y�!B����麙-Xo��XHlC��`T%d$�\P�'0.���l�N�Iȱ��4��x�1�K�����Z~�C�f	�LY�p&[iL�X7�=����Am�+~�s�}�J�y��t�8�c�9��|P�q־�����S���ٔ�ѕ���@�Rh��;Di����e�H"�u��T�E���T��b4������.:���Zv�wXu��@�͗mx*��.���yB$aϟ� ϒ_�"�6+:HB�2ڢ9,q0M40��u�~�,�s��
�=�����"����d@�d:�G-����T�gs��=I��qo���������������p)��ƙ�`m���rX���>P�<�y�h�~O��2�P��K}U�����>?��zǪ�~�Ө������D�I�m����c_ȍ�RXU�7XX�" p��ƻ�7���y4Q��S�&�J�W>}�f�����[�>$l;�i�b�n��tE�!$G !	]hя���aSp�#�$��3Ѕpp��2BMRU��>x+щg@�[���$��[[<��2$dՂ�M��%��f��yYZ-v�/Q���Q��K����B��m�l�e��>�@�$�n��,�џ�[��^}ٶ������_�N�D�Y��e?��d>o}��!o�Qڪ�ni�Cx�ٜ�z��6)���q$���ܟu��>�m�(.�o��q��J�Wn�>�-��ExL�����A� |�p z��~ꕡ��I��%t��;��qokˁ��O�+���%Ǥ���U�N5�@F6���)��}g�+����"N�.��Q�d��?�k�`K�c�wնH�����ƈ�&��c�gw�cR6��_I�U�I�h��!����v�l���O��f�ż���8��]I�Y�#2�kG|q�eB���K�:��=��9`ݿ�����e�K�D
�ڷ����L�`�sê�\�Z���ǲ�t�xx�s����+^���:���8�5� !�1����� I��,j*y���5D'6E�24�\���_��M�rG��Ǯ#�&��{8��,~I�D̶�KC��d�)n�QL�����M�G_�9HN����d3���c�9,��p���6���6�3����$��\���I�l������C���J�F+f�8!��<��ձt�E�"�~^9�m� eȏ��<�E�o�+�n�&&/&%����6�Z�m��',����?�?_�{Q�"���2!�og3�~6��JW-��^\U@��Q���w�h�Ga�z��#��u�6���v��=G��ڞO;<B��.1��Hf��mR)�43T�7�4��'����4f��;ğ�E�@�O��~NSG�r��b��1�q��Y��!����O�3��j��z3wIJ����<��rQFQ�-Cnbv�q�HŦ�9���Z�I�B ٥�Tbp�5K�0hݤ�j�������l�����U�*�GU$�d��N��W�K%�~�X�;I)�Ĝ'h2&UeP�hDhf�o�AKy������Q��l_4�˃|�^Ś�̂� y������g>���3��C@A$_3/:�R���͢tm��Tz��z3�<Tnɛ�[�!Hm��u��Y �Å�M�~���ׂk��k���^a6 ��Ø�šN�]-��Y?.H������W�:����L��
Q��W���::�!v��60V!�.Δ鯙L�ώ���9?�@h'��k�#՝Qf7�}SR�x�sZ�@�Y�i:�q�������̉$���o�u,��@�|�t Uxe�hA^���N�\13�1ya��C��f�F������]X"�`P�,��P@�7�h���pA#�`��:���%t�W͕{
��zǅr@�`;���0�r(_]�U�[�up�F�I��¨������YyK��E���Z߯��+#�U�]R���@�an�SP~�dB��*D�*�󎵷�u���<2������Z��K�ʄ�κ��>��b`�,І�*P�[�;a����=�e���aj�k>}��h6�(4��d��c-"go�O5��U�(<[�+�$�R>��A���>1������WFu���89���v��Y`+L �����9��v����
l�L��BXux�#[�e^}5���u�CZ}�V���6��G	+��kZ�N���p�� aa�&�Tb���������D�����f8���� �����3U�u�smIM��2�+{�u@7�%�!t�K��NH��r8�b����������T_~$BOK����O;RU�G �/$��G=�,NJbW�q]e*����ke�z7����Et�� ��񒳖%�ﭪ]�>�
M^�lnl�������Y	�n�H�_��ꃱ�Y����������@�_����w�.�%+���o����_���L��o��
�̈́p?Zec�C�8h�~�ٛh?��R����?�Έ�1]�R�'�)F��5ol@��)*�ᑺ��R���$�.��>' ��X=��=�b� "}��AY�š��}0�1v=���K�#/���Z����OQ�M@Qf�0S��_ޒ�Q���(#�4�~�4
�ԣ�4�Js7�d�J����:Ŧ5��r,`a�5�hSߧW��}P,�·ge(��Y��c\U�`8����I�㗧��d�BA�乄�=Z�G�8I��A��ߥ*n9o(�MA��+�=�L���g-ϖdk�8�"�~�K}�@xy�b.8�4���Fڰ��3��,����T��7�v������,��)֨�v_�T�as���$Ea�S3'���"�n�/��-�@�?_]�&X���/�G���rmw^x��Z�dvJ��,g
2�3FBd���X�a�KT��S�=�ݙ�@�⺻�� =rtM���m��y�V��R��$�����*R7	�������ʵ,M�f��P|��_���᥽�a�'�D���K���ݝTH�+P�e!��s���^���@}�']R.��V�<��'n��g��������>��٦{>���\����E�)ݬ�Q��Q_��&ݒ��x��S� D��!,ɠq!�w�SP�P�����3Vj�ڙ7�4W�	������,:��f��0�g�P�OY
�6��0(�@bɛ�\mg��e��+=A��^|�P�xpf`\����w�f�/C��ّm|S�=R��^5��/�P�Ѫ ^���A�z\�P>u�:u��Ô��Ǭm>?�����~��d\]�y�u��N5yKԁ�luj�f���쭸"rc��r/�r �SfC���z�3��
�a�&}7H�v���Z�^jq���5N���`��+���6�A���:2��1m�V�$��?�:����G���d����
�Eq�/J��[�ĞC�Ӱ|M%w�l�%?�����,��1j5B����Δa�!ʵ�}�i;�Pq��DWPC��{3V��͟
Q3�&X�xB����aUފ�:8k<K�ק�pX��"#��F�4m�"ǿ���\l*(#��u���}f<5�{3�LY<�f
��_5�_c�/�됼���+�z�23@���Յ��L�&�6E��
�H���	�-���U��@ܟ�ʐ�a+n�<����oS?D�AeԆlN��=c�������>,�%��HTL�6���X���@~6W��k20mzl�~��ڪxn	�����9*Vެ���<=������kO�Sq!�E��E�Ni@a�.�:��cq�G�Ġ�*�fg����v�ڸ+��|�W3$|�'I�;E�զ���5zg2�?0�!�щ�g\t*]�s:�_v .�l%�%Rc�If���B�<�뀇GeR9T�3�e��K0f������R%^Ƨ�(|C�@4_L�p\�h�H�,�r��"q�(H]fܻA�hW�twX��X�]Ѕ �.�<�T��c�Y@X��4�$�7ܪ:�aA�u����r���}��k�����W���\1�����T���ݤ��1Y��U�?)��A=�A���u�a�/`��d��(��aw������oF�7�7�y�X�h���Q��C684&��K�E,�8_klXڇw�&B��b��=�5�M?�@�y���ゆ��,tz3���0o/WP9�����Xk�l���n]"�|�������r	�k�����"VLt����UI�u���$����ݟb �Ԙ��h�2�U��Fw��*�2�.آ�n �.2:W���e�!�R����{ؒb���[2�R��;p�B�ܺ
���p-C���	��*��|7.T��~�rEĕ�k(@������vV�!L2=��IĠV�a�&BU�+�ͶM�c���\�ƣ�r�\%���p��&�Պ"��r���1��avxN/A��^
8�v�����.���_�D����xtQD �B��y�g;}��T�%�Oo�%�4�#*��`{u3)`�|?�oqֆ�
~jX�-M�\8S	&�O\���*n�|T�T�`���^���<�Dbx�Fu�pL30��u*�ý�M��	��1N�����&�B��('>4�����C��Up���@�\��k;$a��@c]}���*�`���.5b�&�iJ��c�6I:e㥘��e��B��P�4m�xA�l!�w�����V1\b�p��JY��[!AϔK�YJ��]\��V
lOAE��j�0K�a?�8��4;���_=]y6�xBx��'��D✒�i��?�ݍ����M�9l3��?�>u�>(FIt}S����'�H:A%�]Z���G�%)zW�j�%bZ��@Q����.��{�����������
�����@���"VJ�G\+⾝]R-���6�C0�
h��f�v3xd94����K�)�H4
�c�\0p[�wYMa��7U�H�H�y���c�~���[%q���RM��l�]#�꽝�P
@0�M�x�EoQr��p�>���:��6�<X��#f�7�(��A����|Z�QF���:͍ư ^�-{�OtJ�"����/���ߕ�=3�?�E5�?A#pQd�>�{
���Ø�&V/���d���zg|����4'
�����['���ȥ��I��RO��Cݰ��m6ߺ3��1�D��^1�v�|V�����c#|0�<�v�������o]H���m���IO��$��G��5>̔\	C�+9��}E��K��&/^5G=V9��ĠT�����k	hIKd�q�Ԉ%r��	n<\�tze&�;��/�V���ݬ�y�Zp����&�Z�9.ᖵg�����j��ɑ%���Eo0�w������*v�Fn��!|Eg�%�fEs	i��S)_F�<�va!)#1H��d��VAW�`#�C%��;��|$L�b��w*[�*��X�__�r4��n3���3H���M{Be�O| e��2�����R\�&k���8c���+�q����:��=	���rK�8T�&[6��ww��B�  ���L��}<	pn�Y���<h���羬���L�zqq�H)�@`����$�:��I�N�Rr�̪j��V{W�Z�TXjJ��C����ϧÅ5L��P?����+
�/1��%m��Jo�0@��v��8" �2�t�*��$�V�0e;38t��?!�w�avL\.�!䗭b���[�:?L���?�UR`�
�̳�Q	��|���&���/����Ůo�������^�1s��j�xgq������[4��Mb(]��AzU��z�k��ȃ���C�,}6����I��k�ubyhO6c@Y@<����r����9�!��ɖ&��G��˒,2YAxͅ v�ן�Á�A{x�O�,�ͣy��k��_����-G�ȟ�3�w'�=�_�]5c#�\���)a4���G�*�b,�(��S0ޜ����qw� |U��:�nmx�dp�{5��(F�N�"�t	<���94�����V���x2�E�0�o�Te4h�)�qf����P���_ѵ::�W	ݴ�	���ӟp5���w˿�h̤f����^b�xۼ�,���߉	F����*T�!<�uo���氨d��E�wl�-^Jv����o�}���oY��Wdc��1�iD杧�=�p���ѳ�љ�X�u{Ӱ{%3���8�b΍kLD���'��-:��d��m�ȶz��P���=��9G������P���m��d��U�
��� �� W��uRn�������m8��P�)_�Q|�To]>EE2����s�R��C���ޞޡ+vB͸����E��$��a��Z�@�d&@O�z(�Lx6�X�Ni�<�uX�5�I�!��T�@�n͐�����
y��1/q�s��蚭)�*�K�K���Q�l�����P&�\��i��!\8iL�ͧX�#ujxNZ`�O�R�U���=/�^wF^ɐ��(9�WI󊼀�k�� >0�C��}o��Cε��k T�u.D��)�{�9���\F�s��ۉ �"F	��ѥR�Pe�m��|+�ŏ̝p�#I��z���r�]%w㔌r��"m�}��a>��b*�O더�.!F:���0?֎�c�³���@!�E0�/Ao^�9��&�	[[��V7�:蔩߄��T=�=�3K��?�2��_ު��Kכp{#E���-kq�T}�.X���`q4�ԝ����.�_8q��[��2�MM�A�@z
�;��q���~{x~O��x�TԜ�=��H����>&�|�G�z ��)f�`I��O�T�8�vI�NOUi�T���1�H~�Ԇ���(x#�Md��1������`]���㼈v O�����=q+k#����I`dv�'Y���
U���®���tvJ̑��_�Hf��xD�� ���ߢ�{�;9����v��a���j�im��Z��у@V�{�R�$U�X*f,�����x�&aK�3]U�"j���x|��x�Aƪ�G;g*�=�9�8~�>���-����%Rs�����~K��{O�ǀ {fӸ$E�*��OhI/9�X�����,mX�F��9��|�<�Xȕ���[��jV����g9��:�"ӟ�Z��S��N�ևk�fu%�[y�v�=@rˉ�,f�����vfN��7�5�On�q�<��F�t8��A�eZ�����'Kp>��k+��3%k�~J)��I�:�K#�;վ^�g��������Y�f�7�o,g:�ϭ��Z0�d	X)����D��^>Dw�O�d��΅���+�<�9' �����\�sA�aڮa�3fQu���s�ɯ��O�g��6y��A���.�{�OrR0I����L�B��^�3!�i�4�3	������A�:��L��4�K8 ���x_�ֶ�d�:��U�n��3�J�%N����%�8�� �Az�{'�òx��ivd半��
�Sm9�}���Цc��?<�����03�]fG<�ij�!���eI����3PK��-mZ��{v��Ok�6�����x쬩.�d�{���F�/SC�ri�Q9}&)�;�����A?֣��]���r�i�+�	���ש���(���Y�.RP��*`��y8���6”�Ks�y|��[�[|���s�3�x'��"d����+�0A�)�kŸ]1��yIgxct���+^���ÓVc��e�D�����W�R~�"y*����]��[���/�7��ny�����pHX���DP���}��[S]��Ŋ�1���{�x)âC�zG��#'l��u:B�~3jSY&�k�r�E
�
c,I�p?S�h�7�+���g�A�ygbq�	s,��Pk��2����4�F��fe��P�N����O2I��S�&u�4s�7����j���I�PC8bR�#�>�����w-�٪}\���#�E�MA��������z�a�XӱG���d'����ecH9��X_�ZD�TŖ��2p��K<�3�m F �c3bG�;Wన׆�4sb�|ii$C�E�����k�Ї��Fy�/|X�GQrW78&�V���84&9(��]V/]^���쀿$��3�0}��M6�U������J
YL8̩>e����W�?�ȷ���wDN�-d�6���b�55W�ϋ ��W�͏lU�%<��)�t�B�^m�W��L�~�����ܳ18��ms+6Js7X��F}����]bڍ����VNҘ�g+K�$P�Q���b�?`�A�r�ֲ�4����
��I:6��)��A����`?�5JIt3�8�J4~�x�M�Ҿ�B~����PΒG�Q�DϞw�k�U�i��V���µW�w�����>ᆥ��kP�B��L�5�:#vf�*���,��3�����k:���O�PSS\���2�O2pgT,.��GK��/�K�
�..iؖ)�16+2<F�\
Tpf���駚Y�r�a�߾�Z����|d� g�׉�G�7(^�S��>�r�tƕ`�$?��pӵ�8�,%��U(����/��uY��Rn�$�4������w}P{�7�H��3�u(0\gZ���
G)��?��/@6c��K���h����]��,�/��]"^O	]E ��Z�r��<��=}(��m�k4կ�	��! ��K���6����r�%��wV+{;]R�V�8�w�W��cjr��Ob�i��CT�ޝh�2�H��rl���l���NӦ�ެͅ���y��|�IC��2��W�*tBuJ������&O�&z��V�-}Aǁ.D����E��B��:����A@�Б�쟀skO�ۏ�gɧE0��+ʌV�9O8��W�o��V)�^-Gh�����`[���R���V��@��kLX�vS�d��KK�"%͑[���>�ᜥ����������'mq��v��}���mśEI+�m�Y�͞��|���'%���DE��g�&z�W��SP;<K鬌L�!SYT4v/�(U�n��X��M0A���+��ȍ�{��p�q\fZ�r1�<��`��U*�B�{p��mo)T2
��u�I�e_AnBk�6i ���Ȳoh5��5�d�l���K��� �y�L�1��y:��+�~i&�W�_:��D�P����6ta&�I!�䜬V��躃��K�4��:�!C>�L6�]���z)�@HjZk��[���"q��������/����Z�L\��R���q?�����2�i	!%����-n��g!~UQ�9b$}~��Y������G��������F�'f��U�rw� Z�@��R ��v�6#��~�>}Q^0�����P\V�����G *��/ W��W쵒?r+V��O��0R�T2J�iW���+x�g�l*��ؖK5�{)�V��,C�O]y�O�Y*Ut��+��һ�������^5g&a�=���>b|7����A��2՞R�~-e���o>�{YR]nT�"�V��ppi�'Kk��(&Vڕx�G7��'^=X@�P�b&?Jպ���-bٯa�b��N��_�����Z���Β�,�H8M�]� #�i��cj��g��:�xz�����	�yY�ܿ�bS�B
0c�vsu��,�~��kS��8�$��1�������Yk��Ҕ_aخ���A��:���[�q^밈�ѱ��r�k�Wy?q� ?>��3�X4M�<��d{~���<]J��VH<e���v�����%��?��	iv�ͳ�d�6���r5���+EI�a�.�5�An���s���uk��w@����6�lm�m��y����Ϳ��iNc0�i]�[���v��藂3�c�i|ɞ� �����mmF�m�FNZ} q���J�L 5~M�;����O�*n������ð>�U�;Ѣ���Sd��P�+��5"�;�p��8�V �GE�ɺ����]c�g�U|p9�@�Ke�QT��xx���4~Y�}�WD�(�!]��?a�����]{s=YzEdң�mnf�3��� ��A���k+zYZ��PG~g?܅�f�e'�X;������0Du�26U�����-����7/�ﴠ���Xj�B^�Q��G���"�K�&�A{|k#�-����h�~��zB.�X��$&�GVfi�P�o<�칸��)��?�+���k��,�R�5:M<q�{?_nՖ��F���B���K��$���N����������Q��ra�A*������4$��3c���F�����DC�����qLzL�b�j��L�=�
bC�n��(��,LY���W����ݥ)�a��(t�N�����bT�OH4P����wÊ+����!ep��ik��"�1����o�[��|��ڕjҸ܎g[�.=^t�K 7Up���]F>Ga�g��#�d��vW�4��y��ot��VZ��H0�}�4��=�Z��I��6�B�ls������7�"�,��
�D�l̑�C�5��3�2���-������$d�1���HbC��GJ��v	 �ra����u�l�_������]-�� �����k�7�zHo��8�p^<�L�o^�\��ɝ��P�$�e�+��xXX���8_��d2��0i���o�����e��t�ft8�n^���K����}�"r�A ��D�d��P�J�R����7"w���3j�	=�R�9�i
\��_`5�*��;��R]T6�,�@�6�j�S��e�+3hH����(,�y�s�u8�ֳCD$,�"_�9y`7M�!��w(o��ᚡ�'��C2`E��=���vv@$�3�_w�eˏM�Y��+���'{s�P�[�o��A]� �&s4��(<���Z���
6�+�C�#DMh������$ŉCN/䜗;�D
�Q���P�GC�z��u�p�[��c*���-�£J���j���:��	St�wp���=S'8�<_��6I���VpuPp}������ؗjH�CI�;&�<�-h��Ҵ݄�;��m�6
+���Hd���@�w��	��<���L��@;0�l���Д��,�GVY�%�7,�1_��_�ҙ��~m�4��5�H�|8���W�ӯ�e�C�:�xEl�v�[���؈e���O�����t*���?��/���藐�i傶F���G)��x7��#�|���~�G8c�
!#�W���;��凯�W{����Ɔ�
-�#��^7�Օ����y/���W��j��T��S��0�$Sa�q$��n�|�D4�j�OЅ�{iy/��i�Yv2�'�b{g_�-6��G��9����r9����A��s8�`����N�nI��k���=��9�
�=�wQ�8J�}�P�P�]B�li*a���z��I���P��k|I�t��3��̈́�]�Cv��}������5��
�r�� %�CO�����<@������������Y5H�o��H�Z#��S�]={=��H��e�ϓ�C`��W��$�&�}�/'>�|Ѝ��w9/��c����K�aO�$	VH g�ǟY�t?�^A�\H�$=�+�Fw�d���)N�9b�%a�)����6 �L����6l�*&I��ѬX)��}���*H:�EL��`ֲ����~}Fq׶bh�}�jCGNo��t!ƍ[���sd�NoH�qTr�b�^G�ay� ���Ə��@GL?��ĭ�_�%�1�>��^���nb��@ɳ� �@4�����3
1��9�K1g��&C�k�lu���hMTg�}m��#�0�ߺ��.N<=�`p8�:B�	��<r�.������n̗����V{h*�x{�����\��ӥ�MX8�L���R��_�ޜ�R5����
ڸ�u=.T���'���e�plB��?D�Й��Bю�H�63�u�X��Դ���H���$��h��6�ZhZ_���Ԓ�����Q�y�w����-1����~Ы��I�5#��5윯9H�n�a+_aD��C�w"a�lHp� ��}���o���<]�>[~;p�/�\�l)菍��k��;����3�u8�QL�	k�d{g�JY�#��.5�<9G.�.�T�'��l��_[���u&�Oy���5��/�Q�!�Q_�{���{s`���̄.G�l2J��^��c�3Y����Y�� dy�n{U��r5��-&(��H�D%�JdT�|��:���z�)̹������/~!j>������wx�?TG��J��ZkY<G�2>�����O��%����!��*���#�!�p�u6�+%�^ ӈ�i��)1Cl���Ez6/*�p7����B�^�����~�$0)�E�:?����V�H���M*#�.�ܫ��^ݞ٧�H�|2t��X�~���Q�=O�t�|w�~V���B'�c,/{��g]�Y���q	��Ta� ���l{B]���D�+����&c��T���ਊ�֍[��hVwp��}	d�NJV�[{T�>Z/�?���gQ.�;�A�6���ɇWt�k�A���XU,�q�ӴbV+�;����Ϣ�\>x��a)��g4�ʋ�IEC���6��$;5	����gt����
�N��Ò"e�F�u��9:l������w֍��G��=�r9Iث�=��	"�%��t�hlTN�P��e�f����d�⩻��aܐ!��.��&Î�X_H�	ː��XO�����Ŋ��TyH��^���/�j�h���+&\5�E�O�#�=������p�Nv�r���+��
$�:��b"2T����g���I)�Z�՞ľ��$���X6��L�WFTS��s����e�O��X^����G��l�ɮr��I_���p�U����̇']�=�I�q4����`a�=�HU�>e�vY�h��/"l����IF��܋�M�"l�����ؙ��z�3] h�j0z�*!la��U�DW�%�a�� ���I��_m8Wm�x����K��,��@(#� WV�^�c Z�찤,��/��.!�쩢���c�8�����w�?�'�,��3�x(``})-l�����)���&DUy �õ}�?#bƺ`}A�x���PM��ȏ� �$u%�f�F��:���h�#�/4�� ��Q��^AA�Y{A�P�߉�8/vfB|_�Z�Y'����x��Eb��]�@�?�	��ʰ ��Ö��#Y�mr����d�Q��V3 ����}���9�$d�R2�D,GH�2��G�a�B��i�X�;�bF���I�m��W���}��!��&�H}��,�Ʉ�������ҩ\l�mr`��&ei8'�7�=A������հ�&����pj+)��Cڻ՞kLޜX���5��0�vp��!�s3�@�4�Mxφ-��
�Ą��;�+�:��f�%,H�K`����[.�[�mf-Q4��ww�^8�sE�\��f�s�L�x�8u�\�
0�M�c�l8
�/�{��[�����qD�,0�8����COϹ-�Y��M{�y٩_����;�H�/���6-�\�k�K��N�YY#k�����Q�Ǖ;;�ȏ�(ꌌ��o�[���e-gK�ۈ����	a��?���-%<U!�Fz��Ј�r@�'��|������̉}��(�����C:�${�����6j�J����	$l��3��`K<G���"A248�gHPR�C�4�@����I�M� ���0,1�de%~���/
����{�b_#f��#��a���ʟ,�y�U��<��@ sý#�S�)6G�K$�s�> n����]J�ľ�Dx��g�Q��;;���¿H���C^�������p\"1�J�>�<(y�F��f�t���>��Ɯ`bT��!8?3.:X���A�s@�ȟ��X���h�Qx�NL�����*Xu=�����+��j����fO'lj��<�$H:�`d�眦9���������"�,]M`i��0�i/ڍ�qe��ǿ:53���xDI]����K�6��ce'[��� �� �GF�~��塉v�s�f��0�Z�6T�t����Zg����-�ů�5V@c�z���KǋZ�I#����;l�d�(׬v��.������?�q6�W=f��U��*gL섀[�y�	p� gDl��<ΛK�F���o��-�q� ������niDȽ��6��?E`I�b�+�]T������6͏ +`b1�^0k��2�%���ٙx����Nf���[�t��N�śWJ���'pdi�j�;�XN;���b@����=�����z)TZH6�Z��c���t��<"�6���&��p�xa U{��g���w�{�eZ�P��~��e��l�e!��.0/'�4k�|=���\B嵴<{�$�@"�����W9$��Ɍ	n��Q����xZ����J��˧���I2+�w/9��3�s64�m��UQ��5���_|����;�9ko<��Xnt%�n'����H�af+SM.Z�Y���L<A�HXh�a�DdUI5�e:�F���7�;脘N��'+�P4T���#i��Z9ng2����X��C)�ĺ����E~i$qh±�*�#5��nz��x��\����+T�X@^��C60�C�a�stk}>��w%��p�h�J^�>������cYQ-�9�;�����'b��$�W���GU���?3�ˍ0*�:k�F-8rVR_Ee�6w���ᙏ4���N%{qaꁍ�Zi2�9�e ��z�ePD�11l��(�""�Z<��NO��.�K��H�P#�M�)��G+Π"��$�S��N��:)CL��
�_ޗ�.��|�z��̜�h�%{EF]a�4#� |����_�o��Y�嗸cL�2�rd�{}�阌>�FZ���`�|�ka�l��{��jἆ�>�Gmoh�G�i�� Q|l\E�HuX�Y4��ܳd�X.B5�gI˨n`�Ƽ��`���Eeɥ%}� h"��Y0[���_띗��\��)<!`Ws����1����g�)<� k�`��Wh���@�B�������'F�;��3�]G11��P�/X�|���ޤ.�M,�3�Z!CG"���?�u����%{��弣��u��K����gM��2�$�G=����nrXu���(G���~�扮cn�Y����}�/--�k�ɜr�P�ֳ� �b�Kޞ������]��*��n8��7)�8KY�2��gA���� W Ŧ�aU����W�/�V���N�y�����}1P� ��Z�>�!�o������I殫�70!�N�W���sw��p2Џ&����{�<��'6>"�C5�~X7FP�{�"��s���*|��ZQ�w�J�h����45;T��M��3��-�����?
Ѻ�M=_SVd����O���U"��V!��#e���X�����U�yU8�H��/H�J(�����$�~����ۮ, J��IC�4}�w�2��lU�f^�bF��9����)�� 9i/:	�9�!��G�Nk������E$�mw���.u#��s�������U�Ɔ4�Op��3��
O}��^���jP	��G@a�3����~��?a�1�-��>���[i�	e�*a�0��}F]ˇ���5�S���N��ò����o-ÈBn�SKm�[�������T��j�ʀ���πO|����Uo�W�Y�J3��|w��S����e��/�_�>(Z`!|K����sbi���n>ԡ"�� Lؘ*9�Ǯ���]�����*z���"�y�QN���@Tx�k�O�$��DL
T�@c}h|�{�X�	Y���KR�'yLϧ���2a�#D��cevn�n4��s��Ҩ�R�R{�9w���t?b|��˭|:M ���Kѻ9`��qi.�\���^#�d��Q����s�IAy�IQ�S�5�i�C*�"�H�^P�i���c0��?l�I
{
� W�RGh?�DJ㬶 �,/3�Iu��L���G��y�l��]8���)4�t��6qf�#���H��$Edo}�|�[��Ft�K�؍�N����≙��#���ja�x����@r��h�=]�WG�
%)�f��I6��9�~P+��fz�Q�r닢D�ki���z[�fb\��~1B��Q�\9��8�ay.)Y3S5�t�ˑ)��D�+M�e;&�U�~ނ�_;'��C��qJ\��B�{�4�0���s_�UH�IKU�f>��	J$�Qx���� �yP4���;���I�(q(s�
u�L�2?�W��p4	��9�Mvfzz��3^�}ֆ�4Jd�FnR�A����!Ԉ�4M�<���~ !�F���0,0$bk����-�iI��K�b$:�+z����T��6w���,l4s�����4FQ+u;��S�Z�#��6��BIׅ��+�ӻE���r_J_�iy��]c��Z�����{,.2����#,1l`�˩B���5�%��(�^�}{���e��.�L��E<wŤ �@Uo�+�a�V���U�6���P�'HU.s�G�������Z:�sy�̙��]��s��,���`�f��8l��B�2g������닩��%헿�E#�����'&T�w�/�~�ƩF�}�N�> 
6!?��o:`|8��ؖ⨯��ڑ"QoqB�6gU�c�����.ܽ�!�.r���䉞^r���G�+�d�nGڄ]*[�h���1��\�7�6�|��ӥ���ذ�V/�Gk0_�Y���-��y�dԺd�Ҟ����1�bF��+j�w7���ٯwHq�A���"^-�X!.=�<���h�	DS\�;�H�W������Q��X��}��#\_[�B�$����6%�M�Z��|n��CkΛG�}W>����f�ڐ�-�Ҡ���3L�-��}�����gٺ�6����!��670�
t:�`7|�dk���a�*:�/nw]O5j4��j���.��T%�eK�}>��"b\���}�}�%���b�,�Dl��h��ٗO��Q�p���5^4PS�.m��[��@a��m���/��-�zo��3R�-0!�	%���X1�o�ق*e�A9�0�Z��~wui�}���6P�V{��{��99C������j�C6�Έ�2�� ˒��lQS��.�0q�Q��a����@�F�ׯ�w<KrW��<7uI��sN0�H�
�~��oա����[�����g�����i�n]��q�����6qoG�.�����o���@��-/�cA���{�����x�o�F�!�<����z�Cu2&���]�3w�V�9�K'C�����m�(�G4�c��+���n@Wk�;Ҹx��]Ζ_u�� =�O��"~�i��X��vP8q�����h��dA�,	�;m`p��Hz��t�U�XT�g�`�{�W�I�8�|�L��}z�t����O&�-kԗǱ�А���
�����=~eOMv�W�ϐa8W���0	nL-B2+l0 ��A���)�U�=蒩�}^�L��9��vHk8�#U)y�
X-��R��0@��2+d�ͳv&?��#&�v��pٛ��6w#Y��ʟ@��{�2���KD|��wk���>~�Ss5Z�/Kʘ��3����Lk��b��)����w�������jy^���*�@U���J�#v��%���Y�=�	�����;��f�z�Y!�������ԴwZ��@�� ~�W;��X����Qn8 e��N(�&9���T�,Tv�t�s��$=���9R�j��KKw;l�AZ�4�2�{�#�.�*��	�PA����w&I�˹�8y��AǊ�[>�k�]/�?֚�������j�g�˕���ɕy���������r��v��T���M5�*�%f�lT߶R�����A!�.ޔ��UT���-��Q���ֵ`�k��,��_�0X�xX����� Um���n�������ǐ��-��5n����T O���$I�CPGXr���$<��ζe���(�C*>���K�OXH� � >���}�v�Y�M�h�F�����H�ז�ǯ����+�p}����r)��0,�/q��vl�$�&��c��A^V`U��S*
�_��O�Uܧ��b�M�`��f��h���"���YCۖz�I3�~{m�
:Ў_?���-�M駏�=��m]�a�2���Y�%-��g�{�7�p�L錜�E6�ę������U��;�u��BO&$G�Nb�Y�^O��{B����uk	W��3B�����w��@�]����ƞ�r@���9~.�+G��Is�ko���W`N�y��"��D�%�Ӧ�@�y�̙IX�*/$�
�lNPA���A��!c�-31� -i\ﱹkL#q8��Ҷ��:�/>�O����bQ5y@4�c�-b�#}c�ǝ���h�i�Ɓu�XW�G��O�q~���kt��CB����:$m�>d{L�#��­�q��nUV{�^��5��v��p��i��|�j/��U�>��?#^��po�|�B׶/��*��'dZ�%y� 6��]�)�%�;_k�X��3=���|6��eͼp���/=�
��� �ᄀz�=���wOnk�����|��b�#,�j��+�X�v��r�!��.xe�i4@�j|��3۲K�Å4�����^&U8U��u�8V��g/�����0}ո��9�CS�p";����?�bK�B��ig��}K�U��z>�5�qܝ�G21E+�Mj��C�Ԋ+��R*k��O��OzپA�C
�z��~��5�
W���$x��V#MXo/��el��g��ݣYQ�C���Ap�N<�XaA5��e�td���[%"� R!�?ql�,ݨ]�����U��+G�����	�C��Dp�X�V3�е]���Z-���\��'�O`����ϓ��ݻ�YN���҇�Al��Q�;����욪��������h���X�+��H�L0�=�X��uL��SW ���돐Ws}W���z��%�CΞ3[�,��ܒ0������c0HRv6���*��K�N�ÒR2R�6�J��hܪ�D/?� qm��G�>��(�Α���_� �l�3u���ΗB)XqcQ�p�-��K�a��sE��g�$"M��1���?���NHEԊڳ�7V6�w��gD��Ê&_�u`��I75j7����H�:�n#���f���8� �$�t ��[n��{c1h�C�Y {A�I(~,��b��x����}:X+��`�i%�7\�����g-Z94Y�h�`���!�8�-w��vo$�>b+�N;f�a���i�c#�9�VN�B+�rXӣ���ܬ.M,ݼ��cZ����Q*���*���@���*�G='uȸ���_Y��@�4~��wՑ�4��\������de�cT���>��$tgF�C�"�@+��ykg n��L��ә(V�8���'�C���B��j���jr[0�)����b�	��Y�5��	�D,"jYh�+���w2�	`�X��㏾�s\le�WY5�?�I���G{�T�;c�'��
�sW��q��EE�!q�������%C���d���&�,�4Rb�d���l�,~���@�r��W�N�fM��Ё,#�@�F��FN�<�~m�&�9D�������/W�C��t����9��x�[���g�����"�R��Fܥ���N�[� q���Юp�E:U�x��Q�{h|/�߃��@�@�Ü���P��ʲ)B��;�/���XR��=�_�$��@���=$�) �R�������9%�������lN��5D�R +Q���4�l�)�����;h�\��0����[;U�z��?9����ם5YܓY��.<�sؙ`Aܘ��i�+?����9�G�#C9���w��\�؍�����:0K[�`4�����Q٘�P�q�����9,�σP���N�et=ѧ���*���N6Z*jc��牏��(O='Bͳ���7����Y�M}�R	e \��X!d��J���w�?WfW��X���%�w;���u��$��=X�:jWU�]ɸ)�A�� �G���F�P��6,�]��{ZH.S.�Ԝ��kv$o3��%l\�E���~���Cф�8PY��H/�iʪ������Zܘ]��=Ty����Y1����uڹ7�C�
�]O������R
�L��٪�H��qbƽ{�V�Z�*c������^�
,yٰ�ke�1����E]N2l~�*zc���t�g+�ھ��rxԧ�2}���(8����)U
.Q�*@/}�`�����e��ׁ���Al3�l���,G��	������Vlx_��*L�����"���@�Ո����7I�=�>~qMr�fE�.�w�ԥ=y_?�+ga/QzZˡ63�b����j�V̛^@⭃N&6]y�,6#��~�R�h�1���Gr|5ĥ,�5��/=o(hdd+���u���?t�Dx��_
�堰=�a������[�/����f�8N�S7$ӞU����Ϻء���O�����R)
h�C��Z����.�W�K�� z*o��F�W?���ߋE����C{�����M��N�wN0�Ӳ�n��@�6�ֿ�Ru0�ٿ��G��W����F���`0 �~sp�2E8J�D�'B�}8����MB�]*Y�k���Pz�k��� >�Q���ThLǾ��rV���P���ي��*��Y��a�O�� ['�KӁe�!wF�޲�{���♰��R����|����� v�n�_t�sl�Zq�[�a�]MEf�V�%P���PDT�E��x�y�[-{���&yO<RE"���>��M�?���\M�U�5J�W�Zۊs�������v������ӭ���ibT�������5�Ʋ퐨_�;�K��V��ob���k��}/�G��x���:�1{�_���N��HΛ��sj$�>+4��^� Y*p�l�U�3���ħi&�4%�Ԋ2ÿ(J��Tε���,�kt����O�G���?���Z��
������� �~�l�i�9��p�^ڬg�Z�y8*i�O�c��lNT|.Ə��g6����Y'�R8�0L_յ҈�,�_'�����&�H��Q�r%ot�?��5�fv3 ��:+j�����)�k�2PjpHr�c���"���aZ�^�iA��
��&C��T�"{��QY`��T:
���V������&JE���#�m�  ��}�^5"��
�i����"�r`���3�v��X�a5���}8a�70c��%���1�Q���&_+h���c�X��i��md�yQH	E[��j���7ǯ[��̾�4~�hc�Rɝνw5n���|�!F{��6_��J?��ހvk����5ƋL=��U� ��ظ��ca��q���80���Y-c�G�:E�_��2�������r-�P�7�����Z~� F8�Js�1rp�uu6(�(m]�i�"-�2�GAo|"@�Ɍ���nq�V&�5���'�f�>o�b���q��`�������JΕaF�4S;w�i���2Q/����J�"B�"�.��A�xYn+�$D,�K��k���^xE�� ���&��(2BN��1g#ְ��L-�)Ѿ�\Mݯ�S#�l�أb���⌷�����3��j[�K�[�s�O�U+�T�����>�͊�e9�`�&��d=?a��m�k~��1Td3q�������Ҝ{bÑ��������lb�&v,Ɵp�W�j��x䲃�x�s��Oj���y�����[�]�XQ���/�نf�N�O����7�Fb�o[ָI�sO��[�h*M�C	�%~�)�~����ə��H�e�����Џ�v�]U~���	5$���#�,N+3�D��f�=����R-&.P��@�J�F��mqD*u�s�5�����G�ykg��� f���e��ڍ�:�Ӈ���1�|���5<j7�m@K3ϡ����I�!p�=.��@��ItF&FCi#�^���"Z�5»~��04�$IJ��&+}+�԰=x�9����a�U����X
p��늲��m	k�HnnŉƷ;��xH��G��UWua^\j�C=���9v��S�b�+z}�9��f��T�dKI��$3���-��[K?�!vxg�J���������J!HCFrR�W��cK@ ���lCZ���DG����^jΉ�U������z����u �M�W�M��9�j{0�1)Ή,S��2I�����^�Z��̸�aN��Ά�uw8�[�?����,rR�ߺ7Vp�x��p�g���\� ����
��d���c���;I+�oZ��M����G��a���/o�k�nM� �<��zR�o��s��y��˰�[ ��qǙ���]�ƴP&�I<��V�(/�Z�Nl���ND��^'�b`���%�$>Qq1�^����]�^�]�/�;�TW{�xEzQ6���Y3n��.P�r�0D'��v]Ag�睨�HR{��np��"S|���oր0�+�6{~Y�T��O>����&�xE���R>����wy h���K��
�&.��4��uC�5��!��UD���~JG����?�����
i��=x����z��I�-�G����̂P��@ 2��b�V��i�L�x~F3�e�]����/��^HZP�V�Y��x�́Y��a�����Z�
���Ki�(���:;�~��&DX�e�#P�!>E��A[p�\2��z������.q�>��Jm�b!������I|o����]J1���r`m'd��j��IK&_�V#��Ql�~!b��2�V��V\Y��&6�L0j��,������]"4�+��9����5Z�|>�~�`,N=f�P�B���)�m��p�]�����˽w���-��ܜ~Id*z����eQ��+�N�3���W�k����W�p�ƍ��lǴD�"�O��8�⯧z_�v7�Fa{�Q�K������5�[?-z��[�P��X�j�Cڅ-�n�0'm����;�X��Ǚ��B��<w�I	�uIZ}ׂ�^-Dj�������5+E���^�n�DV���>T$`fX=1{&g�2	Z��N;�x��q�>�#!-heԚ��&rJn ���!�K_���3
N�?��M\)8�]�n����9�D���5��*-j;&|W���;����%�����:`b��[���O�ę��\։+��-d����eH)�A�Qtp�����9H���^��<��K�qz��R�����|��[�rc;-��y~ո7�z/�mB��M�vV���TU�+��-�yo�3t]Y�@�!HY^�X�$ۂ4�F�9�5�r�'5u8���qښ)��A�"}�Tσ�2�z��lв%���O�Ò3��.��;���>����@����?,���O�+|�cu�|G^����KQ��f7�<����d�/�����z�ʞh���1g�h�ٸU�m�#���1^������3�Hl;�*�������Ku��',�)
���1V��)AG��R_�S��@"�u�W��vQ����N��Wo(����Z�I�:<�M=g�f,c��D͖?=-������!n��N�������HF6Ϻ=f�\%�)��䫣	/L</C�L�{m0�u]�m��\e��+�'4�X�}��`�;N����*������%���.E���^67ĥ��^ӣ�A��d�a߉2%�Z�O���+���y_Nq1t���9���^ښQ�j�<�v�Z��-�����8%�����_i�G?s�Y�D�;';�{`�k(�w����;ř��)�ڣe�LKyC���վͧ{���O�����d����}��2h�OC�$��5��������r`b�(��e��g�\V��yn�|+
y�� ��Zo�¤���-W�\yBl`�ijL́�|"gb (0!%G~��H2o���XgD/��M��&��p�`{?� �SN!����=�K�
«ڭ���5�����DM`ءGۥ�n<Wo�:�3�>��.��΃�д���7f������J��s��Ygx)6��+���_b2�q�m�e@�wTwq�����b{Y���f,�3���2z$�u���Ak��f"`��E4��Z3�f��ԺG;H��]��S~��u��%p�;I���_(���?D��eQHX,�0�8u;��wb�s��I.�Oࡷ^��H6�L)�h�P0'��}X䪉���؎O��u�����3����ͩ��[ĵf{�͉�k���"���oC竴��r� �� *e8��U�;�W䷼���oE��g�X}zmW�5����+z��9čwvT����o�>7"N[Pȱ {����]h�u��ʪ�M��NGP���5�C1��"�^&��F�E��6�#vՌ�	���Ƿu@�ˉo��N��7�)��/uzS˝��K�ge$䮁�0*���Y\��е���\�PR�z	F��6��ʖKe���80�(Xu����&�uI���6��7�֐�d^ M�0�?���ݠ/k^J�Ʌ�����,��50�3�^��{�������������1rO �w��N���ߙ�/~8h�́T@Z|c���+��0��rv�3)�\�cP��[R����!r�K�T�2&�j�DڶC20�Ο�rg�I:7���r��3����H��L�����::⹈ނ�M��X�=��qCk���Y���	�ͷ�ڋ?j��9�y�@]�6��vP��Z���u�Z@�9��2)�g-�Pc����ֶy�Ί�2�-���!�o���9Jߜ��l8}Y�ZSK���f����C�=$Tބ��.r���RV�Z�cT�vM2�_�e�Rع���da��$�>J���ߢ�w��� ��!]VCy ~����cҼg���u=�]��&_{��f:��U�V�s|�	���Z��X���b�^.A�ΈL�y�^�R����/&���=J��xg��{����� ����  d *��̉�A��!ᛳ�3L8�
/���Q8��V��E�A���g�*��p���`jm����3����� K�0zp*���1��^t�X�����#��Йl|���6c yNk���~ ���_��{�5��;%����Mtu9�J"���F�f�g#�c��ȓ���t��F�����&�hd����r�$�}[�f`z��7�Cc5r���&@��J�P�58+�[a2���:��Z��ԋ�)<g�PB����@�R�{v��7 ��a���)�c��)<�*����F^�v�r5����~�����t�1s0����q4�Z��e���ƭ,�I��a�ǃx�$���l�@�+T֡*�n��'}#Ie�cR��7Wd �������V���h)�\6Y��o/'"�'�٧muGht�l#��wk{Ҁ���txg���
��@�]C��~�.��0�A�w�Uj����EA�&>�xs�=�r��;�Z�f�u���T��Ƥ��{W��#^�٤Y��&������#}��#��i 5�/<%�� ��.J"
�8������dkY2�P[ �#�E���e��T��~���!-2î, 7�(��OC�Z�kZ�_P�
J7���r ��cC` �c�|J��+P =�Q4��J��< ���K�O�^z���:�ʋ����aLG�f-��i�Gq�֡�����@�j���h}o�py�J3$��YHvY_�L�v���͇��MOVHº-��߫�+�|�	��`�@ikh�f�����GB��d���5Y'���� ��0��}?��&�j)��Iis��i�.E?;!j�Mk9N�5
�C_
sH��#������3����"o6K��O��٫�eo�&eyVkP81�X�����8�� ;�W���h��]!�߁���$Н��'=gٔ���Pw
=yV��~+��ʰ
ӕ�c1�Q0ˁ�%&��˭��:���1�ڕӲZvbiwZ�S�uIB߄1'�B`������������<�Y����_��s��Xʀ�TPr�u�mk�a�g}�aE]K�1��1hO]壑.fNv²��b��~��3�
L�Z-!��l����_zJ��E�X�Ϣ�+n-(�c2��؀<HP����WO��=��N(�eR,�!��Pca>ǔ@��DBg�gN��m�o*�fBɨS�=n�Y�8�f{�Uep���1u�UaLJ�R/��>���{w��I�u���5;��-�ԁ���i��/�>�͂`ֽ�\��YH��^I~�ZkR������N*^H�{�||�^h�®�A��m\������ue+4�|� �e���A���<�oF7"j'��8?Uʏ�����D�b���������G���9:�*�F����`r0��$.�7o"�B�Y���:��K,',�
�5�s!JXi� ����.*w�u�-��4���Op6���yYLUT�xq�7Oj�:��ԁ�HmF�P�$�k4�)ҁ|�vO]�`��B��Ҿȿ�s�&��h����]������W"b���Jv��F�0^{G����pȬ��@�ǭ 鲛,BOհr拾Pø�2�;5�K�6�|_��Cܦ؝�[�i�ǆ��k{��]�N1��w:��q����e7f��<ߠ�PޙK����@G%98�J��LrU��_)íZ� �����ڴ"	���ecd<��?tӖ4ȅX1HCs��n3Y��＠bS_�[��Mf<t/���B�L�c%�Y���ϩ����ԧn�<{~k3U*��9Īq�`|.jG�z�TH�AZ;&�b{3B[�l�R���ש;���?)�m���N������<������H��k��2$�M�QETr��I)��d<�C�9즀LN%R�x����9 ���,�E��SbhI���W���+�;�5�Öm�ꬼ:�b�����l��F�F\��?9,׬��%�6)5�7qt�QT�?�Eq��MI�ܐ�����g���-FM}�iWa��^�2r�2���.� 1�/�/���M'���J������y��>blT2����`���Z�6Ѳ���/u"�q-�Y��m %�h�IZ��|���.�-z���ː����`�S6����;.6�io��u`%�x�����7�Vr��@������R���[~��e��BG#8�����i�--���R,�n}���˫Q;�=IӉ��?O�>q�6�R�s��.3�:ֲ�>�|��W��4���=�����t�y�P+�=��$~؄��y��¬�d��w����{�%�ʐ�vp�(���M겂OY��5�zZNc��0b%۵�a�w'�;�f7a^�kqc��RK?T2&�\�T1��[:��؁�9���C����/��,����ػ�12����R�WHp�}d���7S#����E��M�ΆP��Π9x�G��'�aoA�G��לt3���E�R6��	G�g:b �~5�Q�����.�=l[^��:T����S���[G�I?e��D�7��Ѡ���1��ߺ+���h�Q�y��X��YZ�e�^�B��9g��:��E�.u�9ʜ���qL���V2��<M���/�ٳ���g[�F��4�4��+�����E��Ǥ�'I��X��V�c�|��g����?q�ȚjC"�Hw?��l)�Id�A�<�יk㤯���|��!i�9�DӐ2�^��a.>�f<T=�����D��}c�,�� �o�u����~93꿧�r,��en�p�!.Z���M����\���IB�T_�6zd��ub��8N�?k��2��A��;�#�\a�Ͼ�ΊM�2��t��n���,�+x$�(�a��u�x��)�!�s�c@T*�^�,]&�!������o��I�9����=y��TS�<r�ƴ�q1,ﶈ�L4qL֡�L�x�� d �ܡs��q}�~���ܠ�]�ݿ3�MR'��}�k
~�5���'����z��1��9��r����� B��*�ɣ<f�pt��2���B��Dg��s��1�!�o��W�}ғD�m��h��Ç)A�����[ڛaH&R�5���3�����*��`�e��Dׇ���f� P<#)Qr&��y؎Q��������iKg�Ga�$��I$��
�RS�(��B:��~���z	=���r�\��i����B~�����s�ۥ����[�j�q�E��������c��e�v��A>�ܝ.�9 Ի!|�5��M�u�L�@$:���$�~5%�P��a,%�諆L�_U��&�J�E^V�q��w�h�b���!�䰘S��lL�]"|��{qÐ�V�1�+q�jƭ;��x���V����$ ���(��=���tH�t;�>��ɢ��.k"1C��0���k�x)_0���V�
B1o���b�����Ӿ�`��"���1mb[�!sprW6mLT�t/㷴)�a<H%FL���W=M��{�I
�J
)oj�s_�׹
���+OΕ;�������4�Qd�J�����H��>u���z�`�F�B@��2�>\
�Ih� ;΍:xb�ս%�W��ȇa�]e[ ù%��>��k��c��&0ps�r�Z�R�苯�@�$��<��-3R8ǖ�u-��R����N�u�Ѷ�'�Q\	�6u7�����\w�t�u�_��SJN�C [�&�#�b��n�}!׵���_�j��!�#dE�T���9H��AD�Q�h�)����Aw�88�z�GW]�Գh�?LZo����[o��sbgjD������<���+�g�����}-��ۉ�����R80�tG�
�#��O����Y	�.�(���9����5d�� ���8��kź�\��p�U��o��qg5�� ;x�A�A-���~U�=o�(t]9ϵ�*��\jB[`
�Q�)���(g���]�6�������]Y�YþT��6����/@]���4�/�HS��1n;�M�һH�i���G�׹y����:���KL��d�p(AW�&"Oݳ���{\�����t���Yǋˍ���[n�9�l��g2�)���k�#Ͽ^�NE�77�_�) �
��	J�=���m�d��p��%����u�����ekl�������?��.�T���D��P��E����2e�8����̳1��_a� I�?Xש��J��?O���		S��""��>��wv��C �-.���~����1\ HLZޏ=z���wH���=yƨ9�ֺ$B�b�jצ������lp
è���o;h���ʕ�t��H�ԇ�|�tn[_����(Ǒ��HjHpz C��@�(r�o2ޝ��������gG�R�/R���R������D��O�U/d�|'�D���u.v���|�Uat��X�TF__�Sd��F�X���e�B�x1�d9m3��r�x����U1]xffIխ=(B�� b1�1+*��M bo�3���"�~E�q\�mlUu��u���]�����Ǜ��!L�d�[j�PO�E�^��ۄ� �$]����S�>��XA��,��.��S��OQԙ��
:�OSm���;Brf�R����I�������ʥ����0� |ښ���%�k����#�:�9�3�)��h�BH�V?�e��t�6���^���O�c��b&�eõ�Q?�2�����z�����ʛ����4^���QD�{оy��W��,<�g7���4Qx>��
��nxn�q��VU����� h�Qn-��]�+� ưʸ�������Yl� �b��	�S���ۜ��9ǋX�{�Un  -�ӳ^�O������8x����y���꽂�&n�ߢ�m;�X�	�������7���g[kM��T�����^��0s��_z��!�/�t{�����g�DQ`��'|}�*���t|��r�C����:�cBro�H�t�{�����JEb�h:����*���״'���gM��Y�߄%1ߥ��� ?�������jզ�B����v��A+k���bB`6��;,�U��?�i�(x�B���9Q�vu�R�×�>���{� ����1k�����P��W�-�PN$*��Cڟ@��}W|iZ��z��De%p}3xZ�kM*^�������AsR�[�E���-1��� C2*�X���8ɾ����{2�i���of<*$��)ih�_�:pr���߶����f�j\�FW"�k��[��<W�����Â�e�7�x��'��&�}���bO��I�a|������]�>�IR-t.^��)��l%���g9G�9��'x�8R�F�*y:(��KX��l���>g^5i������X�Rd������,g���E2>�?|z�4(}	L���F�2#��_'!�~��yO@�P]Ʒ�v�Z�<ܺCU���w$�3�=b%��6\N4'X���;m���gO4G��.�_I)�zB9����!a"�����$�SCU/ [%|�)D��F��=��΄������9��U��v���{<(���%�US쏆ˌS�	(:�����kj6�[ i>+�g/]\w�s���|���(]�<q�]�d��"ꢘ�7.���W�Cٰ�So�˕�����	�jv,VR|�Qr�[e6���7?�����_bh���KsqW��9��
�w�{]ΉK��ƕܱ9O�%m�v��ʽ���`�nn�3�����H6}lk�O4f幰|�r��o=���Z �A�����r�u�]��ȱ̈n]=��1o_>���I`.�c�m+�ny@�zme���$��v�$kUga*x�\|꾻��yU����թ /�jb���䊬���g�H���U���F��#�9���EE�:�e+,�w8��}%b���z�6�,�$��@�O��Dv-7Y�A���7V��V�0 ۵�~V�����k)r�#�(wa�~���<�}k�s2�(��|�������=U��)l��)E���r����`n��V��IIp{*T6��`>S��'�a��M64��h@f�ڟ"�w.�B2�������E+�g;��lϮ���I�B�;"X��:̴Cv!)�g�Av�Q��b���5BC�oD�7�]��c���qCk�Si9��{���@&ϭ75z/~/�=l?����Uc.U~� �Y_r�a�Z�%�bJ�����Lx�5��F�;8>��N(rRv%@~)/#�rj�(5s}�������SGa۶\�`��x��$<�R�TmK�Q+�6sr�:������H<��t�?cXT���f�����̦���W|��l��ϻ7�\��M(wEU�OSc��]�VJ&BST>!�\�P���f`�syL�����������y�Du
��=)�6�����8y� {�W�}i%*����Z�>�g:-wS��&[���Y����m^+��+9ޭ�vv��r��<*���yयB��/jzt����%i�Zb�h{Q�S��E�x;y���i�(�t(�����<�fH!���3�w�����آ;H�#U��l*�������h�4�f�3W>�lKX�lLzu���a4����	��!3�,"2o��}Q~�F�ݩׅl���J���N�
�d�������N��ѕq��%�����n�
y���VJ����QE�S����`�|��T��J.�-�`�H!^��@��۸�X͉�L�>�+�Q����p�!�/0un�}��C5t��{a���m�����iV���#�;��w?SYɇ�t(%��(/�����;@H�NN�`E6U�?�����!jUw��hԝ�׃qsl��Ԥ��Ƌ�~KZ[�q<E�@�1C�xub���m�ǻ������)�H?�,a����O౎��i8�W�eӓSU����3e9t�ƽ��%���Z�G�W�w���W��Z�.���:��:�#˩���%	�/ؤ�S����~�ͼ4�Gr�J6s�,$m��:5�XB4G`�H��P"R���aNEҧ����=ޛF� %Y���ރ�Lb��l�Q~���m�X2��i���.k�G��!i�Q��7��ʾ��N).K�/T�� CU�aϫ�6ᴮ�uJ~���W%1����J0�������<G|ɷ�mU��~��g�0,��$��El�ӿ�H�%6��8�!��7��昔�
�M{��h��?���z0�;*�F����ùpB*�0�ci<F�l`�Z�Úw���=��h�ۊt��Ć�ݞ�)���:JS�'jN�K?\�>ɐ6^�B���݅�<����.�t�_�u�kn�a���hZ��YnPB���U۞ };�� ���t�k�rϳ�s���h��m+P��U*2��,=��(#����ƫ�#��ݿ��צR�M�/�]o�Y�JY���R��@�n�$*t'��ҽx���\�V���j׆4�����9jWS��7�M����Nbn`_ϗP���1��l������sw&���oi�K��ð�	� ������-���|���J� 4�	��r��v�X�`�ML(����L�y7N)&�A�"4%���m�qq�����螈��qU���Ѻ�.fմ��5n�wr�wF���(��yM�. M�
qe>� 1��>�䁜��)JU�bȡE��!p���6"Yu�_
Ը'�kn�ï��OҤSD�B�sN�l�:�*���O�B���&), !���`��[�ښ��=�W��E.Y^�{l�ѯ�%Jj�^(�}ϡ���p��<c�=MF�k�6;�A]T	y*4����K�y���)Ⱥ��v�:#r ����g~�W,���2?|D��nܹ�2	f���X1&Vݩ��e5���� ����/d�4UX*�bO�����%�w\��,��Vq�Le���6#�Nn��I�$��r�.; �}�J���oc� <�U>gM���ϐ_|_� �Ե��x��,��T�Ϯ�V���H�wM �~�E���lǀ�ӦU,.	"��|{�>P�.LJ��<��2Ǖ'm&B��*�C��|�&��p+{�7�8������%A�")��Id�4�^�7�v��1�]J�\~��ܗu^�n5Q2����e2�c�h�������/â��~嬂tiJ=��}���m�~��xU=����q~A'��{cC��㡓e2�ԟC�s�!.�4�� }�����q3��.���ܝ��5�~�Yh���f#�\��aD���Ә.\�Չj�(��nEY�[�Ǳ��n��kj���Z�d��T��x�O�@ԩ#ǎ8�	j�,��������iZ��5�sH�����=J�X��Q�'ئv�-zA���#�-�	�=��#��?�k�=�nUI:�KpE����h&�� �]W�e���4�Z���;�
J�ރ���f���j�3�d�]G��I�������0CN��@�
� Ŕ�����qtA��~�kZyN�7=e��}L��XZ�F_�lk���mm��wތ7�Xd݅d��������H���J>����+�N]�J���S�7�>�E�Z��̘�����˪�����CD�}�	�.��F57�n�`�v��>`dB9��A��mW�.->\��W�ҌV���"�N��z֞7	fQkO2��i�\�1����D�W�6$S��LsO����qV=�$Q�����A>�F4�������pc� ��?�e���c探�n^���#���ך�C[�%��F5���h���q��ǧ��<��Ƈ�S�j~���-|��&1�i\�5�o���؉�l͞�x�,¼�rf�"�2�m�a�0�c���rT�_�. �
�!����Z��/��%b�0l'0��|�n�5�ۦ�{���@��E���"�ޭ7�m&;�ՙ�p�<s�,|��T����G�m��|-���;Doc͵��A�
e��;K�2xw$����k���<�� ���]��)�p-nJ�J/t�D��'�|� ̸��V�>4�lSU���Sz�jDا	K��
��-v�ň�cs{N6��~�]u�r �l�A5P���8��;\�1Qm��\fc��|���y'���@kϝ�W��-���3�:^����9�'|7EP�Ֆ��­?Q��K��E͆���I$J�/�Q�+����^��E�Z�j�W'9�����6�7�.-Q��A�aby�^	%C��">�v��_+�����I���xz���m0������:����M���V�<9��=i�K���Of�G�F*��õt��&l��0�p��le�*�>�r�@n~���g)�H�����i�hxfIY(���������\��B�;����߿a�EHL�\s�X}���$"7	g��r�!=P��IzlH�^�������F@W��JTM�����A�&bɁ3�eܱ���.XȒp�M�"�n�BB��n~#0����(~�|9T!\xюr�'	Y���r/;;ʸ����f�����smS%���r"C��=�de����x�Ok-0Y�JJuvOp�{���	ĠW%�&�T�~#�ud26��X���+��(0��YM�_�=cN[Z3_���A\�]>>��37������(�������j黈�	��f4;�7Ra��隣H��Ӟ�"��\�J�D^$4��NR����9��^�M5���y�ft��?����c�EO��ȱ��ݒNU�K��y{w�r$�;$����+�K�wO\�:�~�:=����AGYHK?fq	� 'DN�g���Σ��Mu�ݯ3+�e�ra==�*Y�o��7n�r���tD��f0��A�h��3s%R����W��b�{{�x.6U����3��;�;�����R���)k���p�~�������nix�6�f���z5�!�k&� S0�N|��?T@�d��:�30	�O�}D�^v������靊����2���Ōc�5x�ӦCӿho��Ŀb��y�jY���!�bE�:�_g�Om��,��W�窫d����E���79ٰ�l7��:_���$��G�-�n�!aB���8��������'����
zV=���T#Ϗ���D8�1,*�8�休3�L.��Q�0ʓM���J�&!����w�D�����Hs)8/Ý(l���S-h\�Q`X�o���s�St���õ^B���z9Z,�l�+$��t�}Y����ñK������-�lV�o�yЮ��m��v��c]�>�0Ch����I�1x�Y:�%�yԭ�o��Iz�:t��u�(Q��T�VU3J�1W+���\&]����T��PM��8/ �g����&�M��Pn;�Nz,��H'J�<*=_�=�DZ��}�CU���B��S�7W�:`^�r�)וo ���]x�E}�{f������K|��Z�� \��W�j1V �{F{7�G��8���W�<5v�9�␵_=�c(�Wr� ��js{�)����ue��?�İ�^Һ6UUj{�[_]�YI�	eKXنz�wE�j�=���X��pt�şE���F��EńZ(�(Xn�b�7�5OUA�Flq���Yy��V`�B۬�峿�|:��u��+��y���{,�@���b���4����
��o-"�-�|���е��$�������,ϗ���N�͛���N؃d�ӴWe(�ק%�����0�#�����ͳ}�#̰�h�%[�5����SJ���ԉ�� ;|:�a�Hr����{��І�����K5~���
j&"�֡�ԌryHe���՚�WL/�@Je�N/aT��頸��i������ܷ��#�ûЧu��w�'�A��_z�0�-8``��si�ϼ��>�BL(y�}_9â<G[���9��O[�����v��B�NɯKF�l� Х������,����ъ}�n{�E{U/eվ�p�`�լ5������e��bsa3T�UืUCY��7�vC�xC[�X���/����b�{������ ,{��1�S���;�M	G���:��(y�bV3�T�S���=���D�}���e��WSG��t��5�2�mÒѾ�m��E9���-+��E4BeH�0-A��Rg�k�!(j�Z^��BqL2������1<�3�f�ҝ+����=��4o��UWX��&�2~=�T&#�q��ܜMQ�E�0|�bႛ��$6��U.#�n����A���MF��L����\�)v�)���if2���-iw�!,��?�mz��������#%��VS)�#^��?綢܆�_����)��/;��|Jf��r[W��8��rӛpv�����h�rhj��$Y����o����f��q�LZQ��q�6�������B�!z�ܲJ�����0By�ur3��s\||��@C��R�d���xЂ��
��J�,;=1�ʢ�7�Qi3��^��U�+���\��X��wh>��Z����L��y��ѽ�_=�~���A$���p��?��&J�w�KfY���A���kJ<��,�}���V!����a��$w�]��Q����ql���W�s����(��I?���Ls�v�I��p5�����Nό�1e����A[��sS�@9����^�ųʭ��ǐə���������{Q�6������]�{!�����|t�ߘ���UǠ(�����j�����I�"}�+��e-�;�	�����?;���A����aU[�5�'8&���J���f��d�$��%.;�5�9��8���cN!1���U`:�
�'qu��I���`�nR��58�Mo�0W�ǀ�D����ң�Q1{�'��33��^���v#MH�r�i�a��Ø��.�θ=�f��{��%�{"4���~�uk�w~&~���bo�[ˈ6���p�~=�%K����*����,=��"���<��,� �@��Qmr^;��B��4��pAr��Ι���B+�lu?GkN������X��V���V�0��i�l��w�oQ>�zm�����*��w2ԁZ�1:!${a���Oϴ-�\����Œ�A� j�Ķ����w-��Kve(�S���L�����Q"�)���0~� ��AY��n��\���u��}:/Ofo�f?�+��r����%q{�Q0�!��$��T��¹����2rf���f�ȷL� ���[�^.iFc�>W���m���-��H�� W��,�&c��V{z�̻c)�7���,������6N��S����`�UgpY��3�U&��,����PI���`�l�%E��D�j�9�ig���2��z	��P�ĵ��D��*�pp�R-��U�}��`��L��܄�:;�{������|�D�f��,�t�a�Hd��Ұ"�ֳ��}��d3N}��J[�!q�K*��s0(����&�����M�fs��,���Qk�h|Z�\��ώXF|PT���Ƈt�~�
@�Y$�d�_�Z��a�_=�%�'������Y����9V"w�cZ��k�����ߊa�"��@�&`��;����Q/��a�/��|�*��~)���Ώ�����N�Qج��-�\�]ov�%�#��2"�t�ۘ�����F�P=���P��#=B�s�o�9u�'6�]�� �m�r�~�`�90��5S4 ��Km|oa���,)p(d<����7n�?M�7[�>���6���9VbA�\!���HG�.�A�NO˄�C�`���]-���nb�N�IP�P�x�p2ŀF�~�F%�_����o�WNg]��=��%-�}o�!@�i��SX�R¬;>\Y���'�.�� �B�&���Y�Q=��MӠ+i=Wz>���
 �?�=�[!-
&����%m���̇1�ё6�X � j�æP��\H��.l�9�9)-3G��s�������Z��M��� ll�7ݺF���KU����K	�lݙ�x$���_\�0vY�l��tE?�9O���u��ܵ���:	���#�LZ�㢍�$�K��1Q���!o2�<��I�Ҝγ���msI�DI�!Y ��,B���j�7�eC/����B�����:n�U�F	���Ji=��:�"0e!�7ylW-��LV��v�f�Ē����<��Pߌ��&r-�ū�s�ȶx��B�"�����ɘT|:��'�)��f����s!�e0������Ψ4�X�ٷ�����(=Ӎp8��o�p����F#@O!�.ل���Pw�1��5uK�����x5_ˬ��"�XO~9��o'E|;����y@���n�, ةֆ�Q`8���0D�}�6Nk�el���Y��{���a�q�T�I���d���]/���ts?	Hc9�|S��Kl����'3�Ar�3���%�uf0�q�ra?ry��D�����y.�3�cToܞ��o(��$L��}�*���V�y��K��l�X�\�����M+�G��r��|���ٺ��c�\�y44�8c}>�k¼�}��ƾ
�E�����b|ﺈy�����0�$O�X��O�%y<����8Գ7��E��L����f�h�cl(�aD�up�Gj�1���!���P$U���6%�U�|�B��Xߏ�e6|��g��Io/Zq�8S������@y��mP�}^.�5;$�Be���rU��x^�P��Feb��̍�wm *��2���	<�g�{���mD�^�oQ!4x=�~N��ƿ���馷5�>-���C�vxF��ēȧ�q�{�QN
&e�q!�1�x��Ħ���GzJ�7�>�.��c�_Y��e(�A�x��<|�G�IE�I��u.�V���'� ��i*ԡ!��}��l��L�\�4g��3�	�� l�����B���q�h<����ģ�Zh;�\,/��� W_Um%ƀ1@���g�VK��]���(����A��������,�����2�����>`yH���$��YW�S���H���	wn���z#6�����v�Lp7(���ٻUį��[���t�jp�n�λ����ܠN�FL�];%�G\i��as5$�S���O�Wi\�Z%�w�g�����p���}���.���q�o��ۃP�,�����^OGZ���㨁a�S�_DL)�P�5i�aD�QG�+x���Ħd<ϼ�i//��P�\d���I�����Gƿ�G��+F{EC�K�-Y�Pj��*ឫ�DU/���|�k�B���)�+1�OBW�?� ��X9�m�q��aEm�]-ť��yk�C�z�!�Wر|L�Q���B��2�����mN;�=A(�5��V�)��m]�fo����*�Ԩ�]ھ�U�b��.��ky](�a��Ű��e�GĎ6��Ʌ�ռ���C�2P�%	����p�~2}���#�J��(걫�$'D!���2�y�*q�b�=�4S��I� ��r���m����Y�ۢr�բ������c�4�I����a
QQ2깎�/�Il��l�������g�C8"�3�����l��ͮ{�E� ��EJX���jZ/��f>��_�s^�֨H9V!������F��Em�e�L@f���Qp� R���Їj���׏�!7�M�L,��@O�kK��^ $;[�es!nD�@��{Z/�M��E^��qq���O{�]\��0r[���Wh�8�����V
���
�����?$��ጥ�{#�2����8�����Y�&ә�I��cA�͠�	r]��z%A֫H���s�[/��Ƨ�n&al	�M�
���^��U��[�J�/�����e�(G�u蒭z�N�j��	q�98�V@�}k�� Sm5U~_. z����8��J�
��3z���& ���V�"jMu�n�\h�$oj5�K�g�ZW\SH���O`gO�;�[�����4���z��"1	����[~	e��a�jw�6��j�CĹ$������ ai	��׆w�$�T��:r��0�-��R��O�#i�/�)T4-�.j���rDs\�G��NH����F�7_47�7�svWx*�LB���M\�yL��T�e�هT%�B�UX��h�Ĵ�Ψ!�$vޯ$jO�d��HB�0�#1�~P�e�PK*���}չ��P�U�6��&U�ꔾ�@ZIElZ˅�Y72B�����(XVsd�s�\i���o�b�J�p���5!�Vؤg_��A.K�Ϸ:�b$�g�9��<�,��z�D�V�O��&eb@����2h��=�X�jx�N-�N�2��ݪ��'77b��%rluY�ͪ������ߚ�ϑH�zyi]�n�Hyy8r6��n�'��g�������W(�O�m��[�y�@�Y�>w�L-g@Msa}PRH���P�T�% ���"��h�B��']�D�i��(l�H�O%��c಩)0���,I�@L��]���}+�l�X^z&���~3wF�F-�!���y�3��p>�B���fXyU���+%x6nO��	�"��}���~�73`�2/�2�a�x�E�����C���s�ik��o�����}�?��qq(�}�t�f�.	�\5�S�2aa����X��|��Sa ��5Ep����7�_<��>10�^�Z��$oh����bs�ԕǞ����a�iBm��I�����<�QZ8k�L�(�"�/QRk}^P��٭�H���/�/����f�6��Ak̸�
16��jѳ1�
@�:h��w��L;{}GZ�f���"�^���|#�CQ&3�+u���l�$�j�]�V������㝎na�̤�-HF����)�̶��[���XV���^�� �L$�A½D�1l�`�a����p ��O�6z����۫o�L����p�����	���7�*J$��j;\Z�
���*p�NeO,?�ϭ���~�D�ְ�d�YBK_)�%ǚ���J?�T�&��2/�Ô
����X�@wK��'|��,��J��h~r�������C{����Ǉ��t�
^I�q��S�G�wy����iSu0y|��=�#���B���{����R��&����?sA��"tc}O��f����N32�U53񌗁ߦHw��-���dg)��AU�O�*U�Z�̟Pi�D;%�e|-KV��h]��o��3�{�ú�\Kޖ��+�NN֍m2�`�D���X�-�ɸ���6�9�;6�R6P��m����P(��=4]Q�kΊ
��V����$�z�[�ꆯ�`����]�bF�%�^U�v�"n��:*b���-�Q�� ���6�s7R�fT~Vu�\Q���,9��9�-&:0��(k�!�<g��,r46�t���l�g��P���nK?%J"�>uMB5_d�yBl���H����΁���_-HN�Z�b�{�lb�/:dy-��IV�����s] ���wR�F���xF����B�Eby�c�6է�wQ�p}yF�	�h[%G��{����TZI�%qou�}��,���>��*.٫�>Q�_���SS�;�[��"��f���pNXh<3v��H�Р�u|%Mv�����/o�Pz�U����'�lM�O�p�V=q�4���g|������4��®�Y�do皌S��pH���sa]��R ��p�S����t{�����X|催��b�J$k�4mpQ�BsG�������8oqTK�#���Z�k㠘pS���N��+|���[�xR��4�PQfQ+�ga�.�.Y���Nּ�p�T��R�0;3'C����Q�T���� s�I��8�������Ze�d&cN]H�K�ڐ^]`���j�`��UK(.-l�AN�Xh���}8�&~֫@q��zG�ť/���^:�6�G?�[�1�2���zp (�*�E-�H1�g>IY�gN��>4����:��Ao�ƴ��[�r�˛O�.d�n܉��A����'��p�H6=iH��,�^~SR?���˱Qj��4��f��3���ЦJj"�I���N���};'�A�h�y��x�]!��@���S��?/�I�d��p��"%��I�L9�NO���M���a�Ќ�R �ܱ��s�F12q�^�����f׬�������JM"��Y����09��׎�갳I�yc�x���3[3��W�|?��פĸ�9©1�[��5�f��k�Ng�]��w���".4	T�k�{�:3���'��Y潸�37'N���b6�m5 +�B��~����nd�z��}q~~�a��mB�N���Q��H6]7Qdu�B�J�W������F[����J����ӱ=�+L�SӂE��5{�T�Z�e
~_���8��8�xjA�=���}W�
d`m��o+�}.��B��3�Ap��'��'�|�按�~��Ω(�T��ҡ�Z�`S��^%[�.ۅz�$-�C�b'����c�b	�5��M�/�G�m�;yES�\\���3AmU9�QH d��[�Y���yf��5�c����S�m�p��`d�a?$�5��A�塞_�`d%���v����x����m�B���)C�f֛��Ἑ��)t�~.̊��L��w�w�(=��!�.�y�_�������S�Hk�@Q�!sӲ'ӓ�K����w��"b����.��o�M2�߆�Ҍͺ����B#2�Ǥ�U�9*�	�Y�'?��EP�e����w	*Y���S4��}"Λ���vD�L��2�%�&LQʪ��֭��\.��:�?%��G�|˽�V�.]�k뼹V˟n!6�n��/Cw!sg�y,���?�'x,�� ���m�{�{:�:6D�l$B��ub��*�A��4yg�,�cBMA[�I��F�{�R�QS�U*���|=��&Ӈj���m�dI�M��Y(Z�!�''B�E��r���w�A�\X�Ȟ]F�F ��ÐxM��,z����,��Jn�N�"CZ������THK�+;�M�0�8�q�ؖ�ipH��O�d u����yI�G�4�)e9��|�f7����3G�e��#�f���X�$.dŹb��C��t��F����a�%+Q0��[���SJ�����F��b��}f @Sɲ�7\�.6bOu���VkN���f�����t�~ ����Y���� z�5(���"i�"�ڥQ�>_�|����T�����k]"����+����k�%֐d�>�u�Oz�y	�I�u~s�T��! ���n�3�h��]����qiW7�l����!�&�v؀�^.c �і�WOY�����-X���A�Aͯp\!d2�B���	�l<_�𺹽���I�:g2x�*S��$�ߑPgp�a����v?�9���a��$Tm�b�g��o���p�W�"XvLX��ZG��1b����������ʕ+�9�@j[-���Mqua����}h������x�n�����=��z�qYmS��>��}�_+�?��d�4������R���T~~��Z����<�k�ǽ3KE�	��g+��bh�|��Lh�Φ>����Y�k�>��˘�?g�s�G馝����F�5��m�;��z���7az�+-�Gx�ϼ�^�1r0���;�_��Jy֠��6�m6�Α�/AsPڨa���ߍ�1K�50���[aO�����`;y��8���tڬ���z>Dq�Њ�����;.�����`[�Z�c��^�%3�G�鋥Y3��R�G( k���IJ<w��X�݁
g�[ث��5��^@9q��5f�����V�cZV{�hǻ�uXk��rMc�&2oÙn"{�V��F�R9ą�ηU,%�6C*Ka5^����.Zc��֧�l��U������2p����TX\d��\�Ѝ���O���ӳ&;�LM�v8�PB��k�.}�M��a"����\W��L?o�K�O˧i�h�� �
��I:���9�۪jD�n-��m��tN��B���~�ȷ�#U�6ￅ R�����R�%k|	=����aaPk�Z�LEnDґ6��'&w�Kvߛ;k'�r^6V�@ȡw�,�Ę@�h�1�`;
7�;�']Y~�o��v=�{�Q�j�}2L�8^9i	jt���0�/6#kƐ�����4���D�������I�A����g��@ʗ �T�ڸ�@�{^�2��oq`k]�\�����%{O��=q������Vt\l�SjDݯ2a�@�o���3���(t mc�䱭�c�q�20����or�[xhN��AdF�Y_Z�y���GJ��Zb��Xfދ���<^g���o�O�KF�=�9S�ڞ{t�G<z�5:@ro�3�"�*��E�.%��2��ޘ�Q����
�ݞ�U�Z�����H�Z������w��\�JQ��y�?��M[K;������7A�P�J�Y�H���d�����R[�fl�N�DIU�q+GJV����Ȑ������k0o�v�A���sy��-�����R�^;�9ՈT�6�P��Fb���/0���#ʭ�	���r8�'�ӹ�P�y�ə��g(�����Y�٣m���8��¼������G�(C�s��Unɉl�}(𐯲"Z�nh�:'4�������^�mA���N3�����z~������G��1�ę	l���/B�"�MD}M8w	"�0��י�~X"�F��$��uXy�kL�n�@�p�y�"}}�8d����M� �/�4<�m��`�q&AB�zjP'����W5E1^�a��y�
31"���R{,z3N7F�=-u �Gf�_Qí�z���s�����߄��9�>�-��-�l��A�|:J�d���4�>BN�?R�'�Ю�B��C��+���㜈av��t�^��di�����g|z��T	�!�t�ekVU7���V3i����}:i����,v��J\2l��"6+���]�
�\���D!�=ן� xK�
p��%%�M��J�1�Za}�}���B�6y)�M�D�V-jm��TW���x��2��)`4���vK�&)i�z�w���(���j�zQ�$?��ex ���C��%��1�`���Af��4L���IN� �������+p����$��*B-o���a׭�o�:�A��{�K2x��]@�-��%PeS?��`�N7Q�i�H�^S�,QP
�cD�C]�>W�=��e�yp�t|�6!y��7˩
�dѣ�q�t`Y�vZ���Sܘ�T�ۏ��. D�W�����Օ�e����r��4�ͤ�235C�y��u�R��w�}~3�
s�Շ������" j0�T��j�5��:&R�l;B��?���n��ν��2�h%	�4���>��j��J�#��]ZgE��o�x�H��:]W�S��v4�~�ܬp�>���S��KĤI�OTQ�d�k�$+�kӳ~(}?:��k�����GGtJ��'T��B0�G�u�]�ߎٞ+X��J����-T���g>�k^��E�_�=8�V��S8�؞�s��a���H
��!1Ο��Y��D�X;z��[MG)��`eN�]]ᇳ�(SM�����j�/��~�'��E�C�u���4nY-u}�s�[���q��~if/�dޓ�ݘ�~ްcW�ue���-7W��)���N��(�̴O�F�>�-��/"��;r�����Ł���W���=�MkM�Z���Fک˧�ƚV��Q��[���Aɨ9���X�粌�$�ڸO/k{� d��@��d޳��:Fm�(?7Vn���u���o5��zߜ��ߥ�,�lq�F;��`j9���T�+hC�;f%�ZU��o�Rk�	���sh��_�ra/Ol�FL�xۘ�H4���-~���
7�0�s�-�=��W�J��
'�f�9�0K�
�-�nu4ȅ-i���n�����]�y���n��y�mw#��uA`�����i-'����������Ǐ��ly����@6�6���&�98��wL���UyG�h��L��ȗ���\���V��Cѐ;UxѸ��nǼ��|yF�<"~��#��IT���O��[{:���=�0e,ng�TPk�*j��v=�8[����f)����%���9�i�'l�3x1�Q��r]��Ğ� Fߍͺ	����K��vz'�H6d�������<·����� �����n�8��H��x�,EZŌj�A[h>�|�D>�][�tI�IjW��=�Gܿ>QY�J���IMtD��gĢ���_~����u�:��5�!�Ϩ�s72���k��Ҷ�"x�Fa�:���J2�?@�K}$8qB+bQ�$�#�ѫ����� R��&�M��ɚOb)Ϫ2e+EP��t��#�T=�.�b��le��7ޛ����q�-p��ܹ���SlV6R�~��{4yGIC�����Y
���b�j��F��������^l��	�Ԛz� ���A����:y�kJ�����yJԉ�q<gH����-tbGIU��]\-J��M7HO�5L�v5�Y�jis�ڹ���?.��X����|8��?�Ic@�r�>a~���8(�e1wd!���l�L�9#��)nmF+íi)���k*Po%�_�mA��I'!ՀI�&y�X�$8)\�rl�	_��݂_��O�8��ϰ�N`4@����A\���C���l�)�}C���H�� �����rD?r�0n�
�G�DsZy��	�M��h{D�oK֝C&ƒs�n�z�9KH�vcL�MZ�C��~\$Z�3*�K�_���G�@�P�.x���c�b���b^K�/�������w?w�N���F�	m��=&�9P�;`�U��Σm�p��+&v|t���P�4��`�����&�ފ��k��U��T��s�����$טT�L��ux/�Bk_�{���1�l�Q�K,�O/ʺ6�
�����a��ܪ�f���q[�[�<� ��|���+Ns}�������kl_��5�ht�2 �F��j�f��촽��1�r�4a���5d��w��iz�uzY�o�QuY�QǢ^Mz�E��.x����q��0�Ro��Z�P��J���υ��ɴ!���}�a��|
�K��az�P�iw��7Cŵ�vy�����<n!�͋���	`�K�����G�!!0w��T*V��[G�?�;��R����?ʽ�V�����}(ш�E6FoFj! ��A�:�����W]��o���:�A�V��$�6>8mX�^ٓ������ć�|.nM�ڂ�?����5Y� C���泑�z�d�\L��o�!�b��B<D��9�i�Y����@���0�e��(�yg3��h�}y�ve8�?�Qu�d���l�Uz>V`��I���CL�<)���K-~�q�∰Sw5ʧ��L��UqۃX%;��X�#�qq
�a�Ws�"�$��P��^��>M���]+��j!c�)���q�q��n�+�̰�����b͌�mE�+��*��zעk0��2���Bc�S�|�^r�Ġ�j����u�Xf���ԕ�l��}��?���5A3���`�	�=�7ڣ_��A�'�潨+��sb���A�Nz���f�-n�X��I�IK�^���I�o<+�����nN�/u�Yf=%t.���a�..g~=erv)5�㸄͎I-�xY�R%>P[.!#�:e�����#8� h�J��H�40��hO���[�Z U�N�o7j6����y��Dpg��B��k�)A4X eϕ����o3���%�n�ڰ)���ԍ��+�_W�j��`:?K�˳0x�?��d6��:
gZ�,L �����	 2��A8_�% �F��c�n�)VG'+��Z�4���6��@��ǎxR:��D�F?��݅��_��Η@�_�Q��Be�C1��3��d�G��6f�K10�d e<�^C&U��(����Lwr�ї@�E��F��߮���Q�@��
n�+>��M�c]Po�ن<j����b���"#j߄���3Xy1P��983?`�b�/JZ��,jI��N�'˥�rL�!�\dSi�Y������&Eސ����bǋ��d�Wj�[b]Q�ls��Q��=g:�� I+v����~�$�(�d�ߴ�gvˡޝ�V]6���^��X4��s���@{_��1K58�����³;�y\(?�� ��n� ��p��4��yL�/� ]�jzP�b�o��A�T��%��x�4��|�W.z��%0�| �+�T���÷���?:O�|�<�	�쬅L��o��Z�gjM��'Q��X�\�~�蝮N�)��A�Va8�y�<ĻґigiD�Q@�����������(s8�(��$�7��`���*�����XÔ��z��ޅݻ�k;�Lva�p��jP(R8V�V�ovG��j��Ae�K�lG��Ř֐��}%{�<�~�,�~6�,�y�fC�/���?]WhÃ�bN��� ���D N!�y��r��+g|�ܦ?�"@ FlFu)v����Q�<�]��6Top�H>�����������O�#�<�^D�\��l�)��eT�`��A���(� j6�D�ѵ)4� �J�qg�$�?��
�Ze(,�IfL�'i����tԈ�#�Ng�c�l�i�_͋���1{צo��r�0�q�,��:4]si���" ���V6��H���������q+Cg���Ҥ �
nzN�^��ɘk�~Ù2j,[k�{�QA$g��%�NA���}�sm��F^k����c� r1�f�}���2o��+�T�V��EA���n�w��eb��_Q�^|�$p�!7(nB�����&� E�2'wA�ԤM����O�)]�޲�R�V�VI�O��$)����ポ���xIRY`[��%M���p��OW �E�oM�g7�A�t&�.�Ţ�g�JrM��hhh��Oz����괏1��_
�d�ű�"8�9) �X]?a�*��3��:7��]���̍F�I���n%)rp�,` ��dt-��龦��TS��f�u��Scw�C;�: k!n���g�i>��~���[ʎ�"?XT����Ri���#*vZ.�i�Q�~�����G��7a,�kh���d$BM�"d_����޴r��}y?��l�l����^A]�eGn�3/$�.�.���=�*�/fx��֦��P�;���sC;�PN�!�(̰��
�P#G=S?�_��NE�Jyh+p�[қ0j��K6�5Ͱ����_�5�
O��'�OI�B�y0�n�����7�rx����3�Q*S�/VT�����LB���V�:��(veX�:j%Ş��������I�N�
]����TG�c�
��5x�r(���.W}��\�$ᰲ�?�>$�|�V-5�	`�`Rq�������ށ�b*`*�B��a�#��B��C�+c�`��T8i�	��
~�Y�e��b�&%3��7h�,�b��O�:���2Il��-/b.HzL�Q=s����]�\G�p�|�9�w�Y�R���:>�S�hTOV5�f�h,��zz�Y���b�.P� ^�HI�����":�ݦ-A6�$_�����n%{W����T\@�?C1�N�	!r�����n?_%x�$��'޹��1�¨5�(4�-�ήE�h_*�u$S�OAΡ�j��r1Յ���_W�B�4����0�Po���eU�/��uo�`���\g/�g�d�sA��2���ɲMC�O#^>W�֣ք�R���ߗF � }HZ_��������6;H�K �T&t]��:ڈ����m��A��I(��
4T�TMHal����M�Q��73V��GW C1*}b⍼58����I�Z��)���7V�7��7C�M���p�O�Z��6����� �KY0FK��
	�����û�)l�%�&h��jo�����+��(=�����S)����{j'��E}Hj�A�����y��z��cʇ��;��o��o|l�\+{ƴ�E��5U8�pB������˻V�6�����m�oք��}����o�Ua�7BOx��i3e��gwb��J� %c�u��5*Qj�3��ô��yw�
��G�����T}�捺GؿU���!D�/�(5��K(H�IQ��V�]��5�R���:Z0��!hVb[p运?�g���jp;PH��/署�B����Y�V��2�V٫ɭ{�J�V�Y`M�d��D3���<l��J�s�v�^s��x�-:9����������,����}a���|�{���˿��������,UGy�(��_D��b>��T>���R�O�-�l��ھXE�;��@�tt�ƚ 3J�ƨk�	��r�:���5hU��F�0P�;ne�ac�Э�Hx�K��_�a�5hPT�x����h�;e�%��F��D�y��:l,T,�u��B�W
�"�\\����~B ��
��6B8�L(�[+.-mKbw`��Ӣg3�^Jy�:�:�'�u�~�^B�cN���X����`��Ph�d�
�H�"ܯ����c��rZ�Z���I��ƚӓ�EZX��Νؔ�6�𕘜H�6-7z���7Q��aIB�W�O^�[F�������?���D��pV���Cr�'�%1�f����a|e���#�˼b%�ߩ�F�t��v�=�NC^��и۪ a��g�m��U��͐��Zm�p�
ec��R���i���,��xV�3�Q�
��������"TG@T\��i�Ｙ��PZ-m.�B���/�ڧ�tT���i&�^"W��DL:6�/�S���c��})�/���y.]�Y�n*�{}����8a�Jy�#a��g�r���E�v���ҍ��=24�J���YtdȳCeܣƾv8�swt��9=O����x�L�n��{�S�}�3[${�L�t�j/zn���脹�^x����;�v�"��3ͯ0>��hw��g1h�ŭ}gy���j��vĠ���!�/w��/&���I9;��m�q�v'Ӌv@	�I�g���E0�ɡBs:_����t�4=�z<*��8k�,\ݢf�Q>��T��aL�������q���P�C�~J���!$���e��4���Bg�e[����rМ��Ύ�SML��\���V���`�"ɾ5a^��{z`���\���nX9��O��:�n=mmng"���<y�nB**�)�i�-���W�-�/�	��
.9w�(#F,O%s潥���%� <��;�@�
z�֓��g�5b��[Q�v�o�h�-��pd�A��=�W2�x+e
�ګ���Z�R3�l��S1RX��'�`�N�à���q�?�C��GR8 +E �@B�@������HV�2*h���ը�z��o/y����M��4i
I!��H�Ј��r���h'^"���4u_���P��?���6�]��q������F)�q��N��	׼F��8��?�ǋ}��Z5��q�|Ri�٫Я�Z��@}�������m�&�N��s� �}��?os�|�h'$z�y���mi���b�|�Jd�T�,_iA-�T	��/o4��(��?7�< �1ϗ�8_�����wk5V�sB�
��U��ߑ!�ߡ�y̲��~v�S�[��U��>���2.��$w�>u�%�|��nI�J����ݟ�$:N�BUN;��5|ю�t��RT#�\�X�*�y�֏"�2����^�Y�&��F:�z��O�yuKpW�N�

�����lH7I2�&I;`lz�I��b�x\�C�~DHa�U8MUw*~M �i��IVDN9»�z�Sh��v��.֡%��ϧX�3�Rn�ݙ�6 |]؋�W�sk:p�78E���߱���i��Vw��s���?�^�k��P��v����q��1$�D:#~��G�"�8
�9�"K�5J�����	��Z���q/�^��W�aF�v�ے>| ���}�9}�p8zj�qM�V�'��+��PKύ@46��]�3���h��g�.}^�����D�m�����UD�m�'�)Y	���3S�4r�\O��q��ӎޮkg�e}�!u�+��HUF���A��5������Ao���e��V�q��l�K���ܙ��q*���u�lͷ%�0�hFD�	��&�]�{��""lgE��ޕ1@���2؞�E��ʣY��c��HFs��K�m�Pj�3j��W��x,Ap�7]�������_Gݓ ~��_:t�A=o̇�F�-�l�f-ј$��1MZL�ߩ�ޜN"��:��ۖ�.N�N�i�hh���9v4�ڸqm@ ��:���s��2O��5[<���?e��J�>Å#X۞�J�[%Zv���8�Uh#��dW�*��5P��cM���&E*h����*rd���$f����5Bo�Ӣ6��w���Eث�[Lˆ�v���J\��'陟J"b�y���D��S)��9���݅A�m�[�ˌh�5�5�%��l|�aƆ��K -���'��7�tl����,T������<�S_ө��&�S��8lm�,�	f3L�l�|u0�sM���U2ڜ6��l�l9O���  �+H�G�j�P�iꄽVm)�D1fY�v�x�6���oG���)R��k�i�:�`!;�{��g��'ϓ��s���%5˷�S f[U g�H]���Ԃ�)�G����\~r��n�M�1q�/_��_���YXC�f��+m�@�N����]_z��� �b5g�DH�l}E`q[��RxM0WG�Z>ۚ�0�f=v��p�`��M�p8��r��2#���b��삋#PBJ,ԕ#��S�R4ІoWH_��p�k(+��$O��kc�V�P�3�u+BF4�Z����4������i�/�Iphc烕��X:E�H/ؤ�U�t>Pì�x鱶cce���.Ih��5:�Y���'�۫���D�W~�����HǞZ�j"�8�U	W��Μ�O"X��R0����N�մ����'r��.N��8F�UAW������|�2��t���A�58��8�d��L-��;��r�`)�J�?��徴G;�e%�-
��~�%B�axn���}Hd�a����c���AT���QJפ\��y��C�݀�iB�)n�F/�+[�\�����@H��
��`ؕ�H��dg��ш�te�a��B�kܮ�/��P��]������������Cz�򙸖lU>HX��SaC�G0G'�Wm������c�i�Qaz���� ;V��z��:,r�4Y���z��0,->���j�ڭ�M]L����C�U�@o*���k��W�u�xb��aR���{&�(mw�o4�z�c.Ls/ �t!o!8�YSxx
BR���
���)�NOIK۔_�k���e��E9��?u�d��]Z�W&�C_��>{���QкV�&�j���!(s X,���U-ѕ&�.�׉������D�T�wF��ML{5D��@h'T��eCqyh��TVR���� U��*���)wOL�ã��{���&��:�YG��~W��	���ǂ@ZZ�����65F����g�!���^'P�)�ժ�lwΩ�fъ[��4W���,�7TEt�h.�ԫ��sa<5�Z��l��e�9����,�6��TEd�X!sѲ� ��}/�8Z��m�	4tƟ�2"h��d��.�0��\�����.O)QҸ��n`�bQ)�e��ފ���b��-�'��A�v��x��T�m;#����ٸ	
���n"��wѕ�ħ�+�\��=kj�7���K���%��5^�FH�{�z�>I�X�ebh�Ѥ��awE�_9"����-(��*(}��v|"�HLL"�����
�q�v�}�1�[��I\j�6�t`�
}DF�?թ�1����p?8���5AxcfL�Kt��ZY�}D	
���U���/MZ�c6j>_�ea�̡��5�u����Y��s�,��>~U-����7������u�W�%���f�NV���OJ@iˢ"Wc��#@�ݼ�z�)�n�^�8����:�-d��غ���p�(<5���@�����>!��&ڒ�����ULT��;i�b|/����W���`�yOV�COD�:�=(�n1�2�_]�xgT��C�[�ު��eL�{;̀����,�"H���pC6�����b]�{��Ҍq�em�����6��V����В�ǂw�r�L�驓 -Z㕮�o���)9�E��"�+�Dj��H(��qס�
�?��$�
�\ ����E/<x�Ԑo���[N����!��j�uv�;�N�b���Ƙ����{��K�8�t�`��T}Ȥ\r����u�p�!(�L�x:��k��H��h%#5d���e��?��:e��p�����hr�H����V +�s#%3�����k�!��u��	��>W��H};�R�+l;�B��h!��D���i L�񋆬<]����H%�G���alt�n�=6�|\�N����JJ������=J�-�M7�;�Rb��+W��}_*���d�|1l�l��"�g�i�H~hu4� �C�N��eӾ��5�io��f�ce5�Z{B��{-=���:��\>��P��6}�{dn|�S������'��/J����ĝ��E#p�d"��i�J�߱��c�&��2;iT��'{G��n8p Z�l5�b��ς�s��}b���U�����J�+1j[��q��c2J8[���~�e|F�J��Uq��@b����3*j�K�(��6��x�� 0�U�;[�Nc�I�wO��������� R���WS�7d������iy?>���q= �S�r�]F��}�Ŗ�N@�I��`�p��W�2��G44A��I�kڿ6R�A�OX��w��(������0T��_Eа�9q�t�(A\523���-��a��_г� �QO�\�:<�;���ȕ�MA�H�s�F
��O(7��/U�rJ6��v�D��@���@�1K��Y~}�,��!���W���W�qLdĹ�ʪ����u|F��>P��S�J��uzX�"� ޱ�s[�`�_ܐ�L���#�|�K#h(v-�2W��O#Kp5!�u@��,x�'��[��񺏫z�A����� ���m#��?�ڔ��Е��=���o^y�-�}���D��*ͯ��/r�R�ȧ��y��
��$��>��o\K�]��p�[E0��a��]��){ƯC�ȧ"a�4��Iqk�Ǥ�Xr�I����Lm��3 H`��}�Sxg���F�~I�2���ȫS�5�!�t�j� ��8�eDH8 ���\_g���y�z>cN-#໰��=��%X|`�����^��-��Έ��Qh3%~���گ�ň�l��d^D��۲na��FS;f���&3����kRn�IL�4u����h���Q�6C~�A���1w�Y.�(��{vϿ��G��.B��n�(�Z�(m� �A��� ��,4��A	��Z�]�g���bT���=�k�%}��]��ZD�`�uH�|F(��۵�i���,�ٿX�b7*��}T��'�>�/��@]��_�?��eM��(B�RZn���t�[N�/qb�Ȯ�t�⏼�;���d��˹��c��$��eȥ$�|aAX��ن9��zњ�Ia@:���b��P�^S�E�_&���Q�c��:��P]E���ݚ�j��Z��H��uy+���@�s�(E�ǯ2e�7M�b�@F�+E��*v��4c,8���Μ���H��?6��/?�����*��k�����3�)9�A�����H���:�� (�`���k���(���g� �,��&%����Q�/�"�/c��$ �q��'0���G�e�qUD�D>�sW����PE��7)X1
�� =,�[��m獲z��R)Q�a�:([���r��%dL�j�i�T��>^S���}�'V�k�C@8�v&?����&�h�����ڄ{�DC�x)�#�g�9*�!����p��ʘX�7~V���-S�^�'�W6�5�|U��Z��r�X�'|�ob����UE�Y�"c�O�+�B���n��]�����%�N��VE�PX�X�M���T��I|�<\�9���bա�7�(����	; 
��QoձI�7�<ZOau�nQ�l����0u�	3A�
S���u��c��E�I��F��O��X'�qE�G&���Ч)U���e��7f�'źݢ��|�n.�A�����.*���<x��!�撘�2Pu�A�\�>g�e�#�>�v�>6��M�:��+˫��ᦺb�F�������N�ٷU�0��W�zEi��5�0�1t�.���/;���7���L���Ї=[����n�-]q�3��d��V��m�-w�-q�*�J-�%,��&x�l>�Ο6!�\w?8��yy�w�}�>���{����et0i� s���v�3�+�>����R���rt'��>>�՝rw���=�g�r~=3{����rV��;9���cg�]���xl�2���?4��:� �%����p
��W
�������7qd��U���e�7(
X����oo�d>�J�-��"���I0n��!�[�u]4�Ū���c��L�U4��v�C��̶����?S��Tbh�r��_@����/�1�^���Ř�1g~�ĥriF���wPl��Hx(c/U���\�w�X�'P}4R��)F�ܱ�5��3���,��a���k:�N�7��`ЌEM}NC�[q�i5׈��=�v���<�U0o4tW%�~�K�� �ȑ7��,f� ŤQX�d�b�]�T��q@t{���"�c�~=��u��9�ħ��?󡋳����ڻC�e�'���7��ݶ��\wg�S���@���`����ԒN���˧Ԫ\Uv���C�}�5aO��5H��X��+����h�6J8(�8�6���[9h�|W�".��h�Cp�� ���8�uV�Fx����Q�̳�� G��Y~��fŃ;�|�e�M��}�Ո�I��;�1�r��.���� ��3�89�()��[>m��w�1���n9h��V�M�,�����e���������/��v{�����͏�@h��+�x�O�mLa�6������S��@���EH�@c�i�/f_Q��#�v��(_ϝ��
\���<D&���ꓯ�א��@r� *`z�E�f926�Q�{�\���|Ò⻅�'�R6Z�R��4V��+ȅ@���I��t��_����Q14�T9���W�Y���"e	MHbA�6A��4��} 2C��2׹K�C��)J��)�L��U���v�)'��m5{���_��v����Hy�}+F��A�n��{IՅ�X�s���k��Y\�5�����T���'�fԐ�e�o�6��M��5���D׳^+��%����۹ �c��̌?��_���EЙ��6�+��Pdw�m�V5qp�{m��VJ���%����R+�~[��l���߱��K�ׄ�wp��~	\Ci^0�%�\�P�A��g��5n�����גȎ��ʞ,�}����N(Y�AO� �՝|A���2UZ���E���G�R��ڏUknt(�&j�L��:�D��A.ڷ��"^l�߲>�_}�^j7n5�lT"��lXw�)�����v-��O�����~��Y�D�6�>;�wD�f�L4q�a]�
1UFiы`�.�D� �ǧ%�oPѥ'k�x�|���'%�3}8� U�Q�f=AF͗�c�8Ś����`k،��w���:��`T��J��qK4vs�
-	�⑇+�N��6an�~���1�+J�`��0�ۼ�ԥ����e��&����5����"�ڞ^eN�q���	�)��W5���C�ͩ�mN�+r�&�>��r��(5��������bk,H��Jl�֭���kJ�`e���� ^2L�)n�k���� ���8֌6��胷vJ	bo%�_�`Q����'Kw{��M�L�C1�w=�"�DHXۺK��3�y���Q�^!U���:�Խ^q_��:U��W�ӑ��c�A��X،����y91�]�O���Ĺ%*{|�g9������U�`���7{�Y|�	���5\mؽm*Iw�+�ROq��ps=���ҷ�M&�{}����&�D/�������N�Wy-�|њ����	F��@��7�Mg�u�&�.e(��.�b$Ø�We���cˀ�-��#��Uqx%ŉ�e��B��&�H����sv�զ��ғ��-��J�W��ܱ>�4'��>��Ӿ��K}ԏ�9��FvSj���6f�����ȌMSŌ%Fj��N���œ�ܼ�ݝĐ/LH\mK��D[D!l��������&�Ӆ��t?��ށ�"��)J�@L�V�t�Gܰ�7@5���\�����~i�u�7A}5Ű�@��|���L���k�T�Z��:Wj��}��:e���]��Jǒ#O�OgQq�ro!��aN)L5�����7��=����6N,�v�Y�yv��i��@�W����}���4aۖex�dذ�p,Ň�n�V��є��y��b�D �ء��Z����OY�E�}y��ut3F3��n��%O`ǉd�6Q3��:�K�ϲ%�����}�ÛA�f����''O]f��r{��R��'�#rCG7=���<9m�֮�i���kn[����4���)��&4�m�/���>��yG�A��!�B7.�v@��E,�$�DPwZ��xs��29����1�Rօ��՚,��8b�Z�,!6�?��C)�2L@��]�W8��u��^�S�+-��c�G%��WW+j��Te�V�&��6�ڴ��L���Vq�٢&�H�I��Mwx�M 2B`$����a|0��O�(1ܺ��̚h�#��ഠ#��c�&'F�?��_@����3�;��)! ���6���z�zyX��VP0A��H�(K�-j�#	�`��2�H�k@�-c�B&����Y3��[�s��!��]�s���E[���%ϱc����\#�޽@�R��̎��	�g��ފ�Fo���Yb�	�j�J'4����^�Q����l�z�$J�ͨ�]���2���ޖ�΄E"�?w+Y=4��r�n�xT��w�����/�u��H.�/�6�Թ��G��(��E���[OV��c����r;��1�h��ęp��T�H,�O��>u&V�B@��ϔj#�:��Ǚg�}���ˆ��7ew����hNb��H��x1'*�V�Y�؋���Q[	U5v�(��hr�I[_���`CPf�>�3͓�E��+i��H´"�^��sΛpޒ��'��q5��,�A��E-mhm���4ϴ� ��@3-}����F�M��_���T	��S<����h�qP���;� ��=����X	΀_����>z>�2Gձ5�O�"��B��G�>u����T=)�H
��"�U<F�/���?ʸ-�~)ݩ?���	��%��@)hA���I��t���~n�df��LݶgMǑ����jKuu_��Z:�B�Y��sB�$i�E��~=�]�c��j�f�J���uw#�2��Vgq��&���V�y�3��}��˸�@�kA�A��MSI�M���Tba�^4�����D�8���eQ��F�]����-�"5��c�/�eI�e\��{\l?2,����	�fo7v}L�$���7��&Q�)�+_���&=a�ط�[l�,p�G���N��L��_`�3Z�X֩�j*`w���Q�#��ys�)��,���G<gG�V#�O�}]�k<�V�rY��?f3�hd���B/9�:���g������{:o�T� w��o���0��$��8�q{����|�b���C�7+�W��d��Z��t����=�H��m���|<�r[�Oo�5�bSY�T|� RZ�/�w��GX��kM!����9����<gN�iG]��S2�Y�䜌,�m<D�5���☋ ��o��kn�哼!Q��:�k��Z�]7&�,|��>W^��(r��s�B��ŅCƘ�׌��{6@B]Y^,:̋������F'�m�Y�{���x����R�÷�!��I���n
x�0�bH#�M�v337BF%�|`�*�!�t�k��.�h��J��p�_Ǿ�EV$�r1E*�~dL�5�� �'"e �`M�gT�b?B�x<������u��YJ��P֯y�?����\���*�s=��Y�h�ɂ	��J�PQG��ﶞ���I�E�,��A�D�i�l�zq�:n�[ýdi�;1����!|d	Y��.�[lx
�| ����aq�n��u_!�ۍ$<*$m@b�u�,I?>@��Qؼ�2��d�TV �#��u�X�%�"6�Lxx=��o�tҤ+)D@�X�tн���g9r�����0䍎�������Qd�N�gw�s�T�ʄ���=��T����7�כ�U;p��.0����{ܮ����H� �~��]/Upc��+S|=��yGq�	״�;�!�@���X�i*��'��]N�/"����oK%�4�9��,�ۉ�SӔ1��j�k:��b� Ed�p��*����n�m���+��m��[U�';A�:t3SkfBl �)��|�}��JBn+������jR]o�Ɔ��So���Y����!㤑)�,-5�oe��!c�^�Mj�O�NPe�9��*�-�) �&9S�J�$n��#���)��3�?5�!H��sq���S��C����S��o1W�ICl߷�e�'>{X6�۰���e$m�K���g*P�˞���kGN\�o�)�r�w�mP�3R0��dO�\��Ʈ�k�Mħ�IQ��g8 ��fh��-�]���ʩ��%�� ��	���C>� �le�,���@K��t(b��'����g
�Y��>9uS��h֣2�q;kF���R�J�0Z��Z2��?�����=v�b���=@~zO�ӂ�
,/L:��9C�%]��h����<��8<�N�χRB��%�{2.�ʀ��_���}�;:h6(n�db���I���C��O��Y��1��0�W�8!Um�V
#�#��(:��x��.9�Y05�S?�أ	1�����5��ugs&��hĮ���������,$�ez^��e�G	�����þ���r�C!�Tg�&*,q��s`���Re��Y�����&�Y�>bz4�F̃�l�hK�����`���s���\9R"�gO��-���`������ģzh�������J]����!�7*��ki���9�M�����e���	��ޫe���P����GҌo�u/cEeG�a����a|����v³�Z�@т�geeh_y	���e"���ͨ�_P&5��B�pPaa{� }P���T�'�EM6��!��m��%Xĭ��|�&G[r$"'����J)�AD|��5*P&o���䝦=��1E�H_�塱]�<;�:�}a�+��$B,mm#{@����2!yFm�ƙP����K�ښX�?�U
�Š�n-/�>���: v�z�:��Y�3 ��� �K�d�, ��60h�;i1�O�G�|�t�]�^8�b�teHؑl�a΢��]�R�;�؂1l\���������`�IZo�c��=�I4��O�2�G�N�yׅ��C�v��s'��]^5�f;���x. �$��֦�I��>���T! ���u�?%Y�4�T�7�]L��}gZ�si/Q�/�H�-��=��� �^�M�P�a3~+���1{�Շ��5H{%�/����~���c�N=�݇Z���^���;����Q��l�
@6O=�׃�|�U�H�뵟q5̪��w����lh�%�W�iՀ#�����Y�տ�O̻;`����`4���PsƇ����c��@>��CϺw��p��S���K�� �н�M?��������z<p���r7��֣���������x�ř|�Z�;�ۄ�〴)��_�U����|�_Q�`�.6���{�}墿p�a���q���,x�
��E�T��X
�a�'��69��\N���t���\�7�Oe*�h~�^U�e��n�hs@��9& ':��.�'��Vj�)�p��X�E�"��c�U�b���Po�ف��ϳ���Ԉx~��\ȩ����	�/�Bp*8L�^�D�|�waD�~���jn��b!I�m]ԳH�*@ܘ��}���+��fU�KL��eB�e�+0��~�5KIH��ė���90�f��ݯ�1��0�s�� �����i�%� 羠]4�M,�h�܇�'X����xwj	0�ڕ&G��O��#H�%\"���<�m�-��e6��kiũ��k��og��c�;�n���*:<qt�{����LUg�t���<�&w`.�U=�D�7;MU��xjOl�N��[�&�Ď���.�eWn?(:���/�s�T.v�B ��Wqe
�~X�&6�p�HlkRFҼy����Aǽ��o	�ƌ�V�:E\��M�./��x�s��A�'�1�+`�~��&ӪĐ�5r�P�w��
Ҥ�0==��)�z+���ό7��\W�-�15�f�$�O��,�v�DI"���'��Q\;���P}��j�`��]�d�0�Q�F�JS�;69�c����1҆&ȼ�����hڈ)���w`{�(LX?0B�@wF<T����ҎcU�H*ZN���a31؆Wv�w����#��T`%�ƨ�!D� }tD"����@y%41�4�@.a1�vOmx=F��G�l��_�Z+l�P�n�� h#�/��L�l�������SZ#x_έ�Z��\��OKM�LWb��	�*�"���G2�\���/�K����+�
 *��ex�����G�;�I�r �����{�m��`��xj`���~��������4�^�d�S'��g\�5��<`Y�r�m�Q_#�S���A��$�m��n@��͹���I��o��I�%�E�ρ�ށ�xb)w{�;a�X� �Lh�M�q��	@��0%=q����H��ۓ�36(V�q���I^fR�U%ئ�#�%|gzg@d�b�,q�٨ٚ�uzG�7{�Z��a�#�B��P��|���.bl;�ޱw�w��V,1_�)�0U]��(y�8\�D*Υ�,o��)��Q����'�̉*\C_E�9u�,.������Hו��Jk0�|d���MS
ՠX�SN	As�]Dtֽ��A%�L��V�YϷ8��Ujc��U�{#Y�z��
��� �m~�2�Sc�t1��yn��`�����>�"Ŧ��-���B������~��9����3EG� �8oy"�ߍBTe!��a�����	�^����9)�b>�j�-�7o�v3H���6�� @ė�ĕ�j��1������:��A�̥���
7�G�ܦis��u�����Mē��֒4�+��s	�3k��~���
���D��C�q��������hs���p��fq�u�Wbw9�x��E�b�����r�'��6	j<v���X�7�z��zP^.X���T��=H�6����^��'&��To�W����z�Cc�%Ψ~��i�9���FY�G�K�a�v�wGgK}�Q��w�בqp��s�_����r���R��U��<i�t�uϮ��ε�2� �#�lr�_B^��� �`���A�i�ׄ�[�"��c�y81"����#Ɨ�9��x���|-���5�F�x&��0w��R����/JO�/���	UcK����*e��q��
��0y������Պ�q��������u��%�K����(����6/x�7�
D���hG(�,���
}9Q��"f�f� �'��4�qU�wv���^I^��B|w���DEۥ�e�z]�+��~/]�)�K&�Fд�t1���j��RB� Lk��q�O�MF`3��3��򓝫Q�����s�ZK��9qɎ�-v}�ܤ{��
ޫY����)<^��������	����sÂa�q�}��I�|^6��'�B=ͻ���5����{��.�ʀ�������w�K
���:��s��ʆ{�B����`�xàr
KĞFTn�8of�|'3q��'��F�Ƥ�:'�'��B�#�E �&�4�U��do�7̈́
��:�X@��?���ˆ�3i�M�K�sz:���~����9�+�'���B��!";�]��Z=/�ɠ
��4~��r�����E?[k`���v5�X�2��utqhB�r��������}�Q���փ��gH������[�'�)���)�j�_��޸̈́TA����$�1R�&�����j�M��>
�� ���s�MK3�B���Ι��Ĭd�I��ST�_��8n��(M��[����8����l���E�=����ra�Ҷ1.>�>I|���th�筫������Hi)��E\���᱾R��y=��PS7��4�(rS��`� �yXha]JQPDn�W�l_*�U����So3�6��ktlj��MO�-}|jJ}������^6]*��{VF��Wu��k�,�5MjZ�����R�s���~�� Mx�?�:C
Z�hT������9���U[���AQOmjDP�Z���9�1�׶ߠ��t�?�x���mO���<Ƞ�~-5��-3yr�mQ�Q��N�֚dB
�@��Ή�0Ǉ͉�|�d��  �_!�-k�7��i2Z��̞Q�5M����"�W��K,5.b]V�t[ZB=-Zj�sR�'K+y�BK�c|�5�u#��yL���W�Z}�����:� l��b�6E-�X�*���;�Ȅz��@�<���W��� `E)}���"��0%��<A�Y�5����޲k�p�ׯR����n��Q[%��:���¡cu���G��q��� �V���Zl������
3���ia-�J����q���u���������|U܄J6JUO�r�:H����M��>�+���Lq����
��٩ߋ���p��#���8�ͺ��v��]��W��4֍ӓ>�״��*JS������c����g�Jo0�ue� ���E	̗7"��x�!f6.t�I1���T�Bo�+z @Z��8I}L�3O oWt��4~Ǔ�(;(��YRo��v�}{ͳ}�Lo.�<\�\��c�,_)X*-��n\��g/0��0Ɔj;��=��1�?���Վ�������p\YU0�txn��|@�5��Ngw��)�q�q`�e���T@����2
D�������<e�#L�Cdg�o�&}β�C�Ll���B|\�.�ugw���Ր^��X��(�|���|Z�Č�P�Ǭa��ӑ
[�����JΣz+�E6"4��M	<@&�d�)	�?>�e��`�gR���F8�s^z��<(�_u1�Z/e�~C� /|vB�o�	-uF��d|�(��j��m8h�:�#>|�t���/J�]��p��U'���G�$��:����V��t��	F�,�H4��ҍ@�QA�d|BQ8.7�+B�'=�p�a�?��2}gJa%�r�?�ZyY1�8PC��Zۋ�eA�	[$��N]o�Z�Xp��� ����n�pش}�w�8�g��C�v���y�r!��wx����@_͔H��^Onb���k�o��0S'9�.�sf���$�A�b��F����Ę1�9ie6�C�ڞj��ߪ�7b6t���4�8�5o u��,[�ӇZ$󣆂�n������i|���yJOY�6K(�� PH.nAq�03#�����;�*Mj���|���=,��h�ԟ�W@N~D5O�����}�U��!�@/R삷�f� �����b�/tr�:���*{��y9e�������DH*Q{�C�0
&D��b��aY��8a�� bUf2���'%���VN��* ���>^�3M��7�)S�>�fW�gx�̽G���Yܛ?� ��[�-Ū� @zvP�5�ݸQ޾���w������?0n/}
X���GA���� ����A(����&/T�.�y���{4]�?�D����GAi����KIO>�3�1�ˣ��K��<��T:C(���YCIcjQR(pziV6~${�l.���9�=a(�'j�����@�Q�5"�.�����=���.�@,��Z�-d���w%ݺ���o�,�7R�O!Y���6ǀ���ާJ���dB#��휐��Ln�G����K�ط��z�`H�3�;�����I;������3��x�-����!��W�Z��n�$@0�R���u�d4�i�~Z�w���V�Z8�`�C+Y�:�0�3A9}�Ea��{
��	p��h�S%v|͋�k�p��]�?{�������X�mJ�I~0� �a\�.@����p�K�MҺ���V�o��L ��W
fK�6�*�:�0�M�Sy�0�:�މ?蜢�~�/�}�����\��>Dd*To'R�DP���0��ͬ�2��Y���6�T�����}4(˟�-�p�-�K�FH�Ì��m��X����M��R��yj��*���X1�g��b�2�@ ԕ��ؕ����^�%;�	<MQ�w,q�;j���C�%���A�tDˎ�b�4�c�(��8����A��j�Z�/Y(�܏�EҐ^"��{��[,�ƻ	g4|SiU��P������{Z,[�����C���-d?~oV�<k����u�������w(^�\�ܬѽN�m�HR��	�΋�I�Ɨ�9K	<�;���w�x��x K-�W�,Ȣd�/%]��,r�H���P�gB��E��i�2���dA"��$w�j���.���z�
�=< b�'�fF2�������cß��@�<0Ӱ(d�(�Qi�7���FϒGu��eh;�,�1�?��W�]����l?2���h=���9݋,�>Ƈ�t��d-��*R��M�
-|K����T�绳������_�H����VǠ�7��o����.}ꚢ�3R�r�|�({z���!'�*oU�����&�	8q��&��-MOg���>g�ȐQ�h���I��F�CV��Rs��oL��Fkh�L��3�8�,�$�������*���A
2�a�B��#�;K)x�6�?��?@���/rC� ֝����px��~?��h���k�����s���k��?�4�߻���_ �Uڵ�]����މ��	Cj>���'��De�^㖲d��zz�yMmI�Ƞ�)�Om�G�Xڛ`��{x17?����.�����jH�4}�Ή?=���� ��tW ��r���f '>:M�
�/H�k����*2]>��0%MF�̺rn&c*��$C�k`> �������[��]��
�ֽ:*���Sq ��q��]H����-i�Uˋ9x�1�kf����S�IeF�m���>�9
S��֥л�����kV��te#�M�>�˶:��B�>Q$����u�,KkF�[��'�<U���ſ��ٽt�8��m���A���O8mq��'U�ڌ;E�o��n\���`HW�a����^i(�� �4;!�rt�M쫌��$��:(I2�1�ob
!'U���1��Pֹ5	��'��z�4�|�>1�XX8E�a3�N+ ?@n�q��Of�#0%cfp�@����iđ˸�K�A�4�vǨ���}z�l���ƺЖ�qg�:�S�����L )j�#<�M�/L�G�
p�)�\�>\���#�i�T��L�^��������\��pg�g�>c�S�3�y�\_���+��N%Y΋;#���#Q�A/�(��
^��=x��؎��:��I�}����u��1��/��c���~������vv�7�C5mf�7Oݭ�+v���R���ߟ�{ �+N6��8ؑ	����״+=)�{�v����&���ğ����nC�cFH���{��&�BX�J�H!�b�_�.^х����h�H�)��+?��͵���-�6~3����� 
J͂�X�*�9��Y^L�0MY׭fC+z��ET��<}!eL	�C=���Ȼ��!���q���9i��Y�G;Zb��1��y7��Q#	�N5��B
�?(eUN���4�*F<��B5�0�;�]�Bz1��@�m	~E�d{t�/�e�؀�1�o&�	�R3�ll��e2��B�Ⱦ������ۡ$A5mJ%��3�&	Rk�b�&8�r�Z8�`M��X��bڪ[��g�)�A0�<󭝝�5h�A�V��TK}+��+.�w�f��K���"O+�P2�MDF�U�y�)͊��!��`�6aa8z�dkL�;�{�.I!�#�ݓz�	&���/��95)��oA����!|�?--]9��֥�lL(�B�º�)]Ȥ�`�F�7�Xi!fz2���i; �Tu}������wk7%���f���z	0����� ��q��T�تS�%R�CG��;����G�pth�9wDq#�L��?�j��"Gh?��!��'�z�"�Hu�U&���t͖���e%��C�T�7���O�_+.������l'��i��.�c�T2�lt-�k�j`bv:�M��r4�S_�8���R�h��i��%�q�Ľ6�&���J����[���B��ԁ�~���&���h�ͱ[Y��vB�8�r����327�o.�ד�fFCo[N��'�"�S��G�V�-��:��!��r���W��7
��������h����i�4�v�4�
Fb�)z�nՋ�UeNI,�PI��DJ�y�]�,=ḃ�s�^"+C/yR�i>�l��O��t�!�¡X�,�Y
��w�� �!��\�o��?�G���|�O���/�v���}��M�7�F����,�2�}�`sQ��p�.*��K��E�N�A"��gT��mL�u1���`؄�Zb����<�*�iS���k8�/��#��f���/�s%����2)j�vwG<|	{�4L#�H��O/�K�l	lT��a��ht�������2M�-��q�{�^�R=&�2�AH��?f�,��)��Qsֽ��j&6�+��n�%R���˄"���K v:6%"\��os!�����I&�_6����/�^�����A4k��?�W�/���r�P9Kз�)�</��kW*X=���(����ƏLpJ,_gpɾ̡Mq���l���UA*��*��kr
��~�o�L0ޘ�͍�P��:��;��3�I*=�@B��$x{&�m9��a����D]�|�:�c�(:�y9�K۳dH�9��<��~����b��2)��1}d_�I}	&B44]���`ll��^����\R������֖�(��ci��d��ho6�Y@k� ���#�,��jnY m�&Z��0�饻�9�7�z�K6*�`�Ӣ�C喘6��D���z'9U��AЇ7_A�S3�&:���om�tG�<f�8�,��s�`��J�IYn껧����u=���X'�Pge������#��8$)�-�uP��z� W���G��6 �~*SuO �C�����cx��	�)Ec��Lv�e���,N*��\�j2*�A��#�!ա]E���4�c�N/�Z�z���]��F������@���F�]�k�4p��H'о���h��z����&s<��Y�'���LuA���y@k���F[�U�]�-�).��8ۂن'�Hi��ی��):b��=��X���CT����P-s������m��I���-�(+�*�l�oFD���6�KkӀt�B7K�.r]`�xv<�lbL�K-��@i��g#F!w娡!Y���kVe~]53�j���M�s�����A9,�m����L
�nح)�������w$�y���&�ɻ�;k�ȋ �ꑶ�[�JD��<�{>���]�����m���u<8l��/�� �
�lѹ��H���~|� a�w�iɵ	��a��ϼGn
�f�ɔ5(\#~�9��Ehc�,���Տ	.��L.o���,��2��i.���7��
j��`���%Vm#IeS�#�`"P��_a���x�i��A�8q?�춯�l�:W����t��3vkп�RQ;�pB��]^�F�R�[�h?`�C�z��za�y�� �Ҡ��= ��t߮�� a}Ղ��<��uj��f>YdKf%�2�Cu��w�yJ��O�V���E� �ln;�Y��9�B��qS<�ڣ�:���n|���a��.\�˭|��t�9�v���tl�;1�mB)7Sm7w�ˢ���i��|5v��G�7&x����߅�<-��A>�[��s���I�E�oɢx�ƩՈ�(籟�Jπ9:̉#G�U�
��F7��Y��-���� ���v����7��rkdAlf.[��8�[%Pok8�CpT*-�q}���7wf�o��Nߴ�\��{���H1A�x��*}=�ۿ�8���L�a�cG �}?���ɨX�r����M���"����x<�r��d�@|���1��QB����� I���H��m����*��׫�����50�D�u=��8�x>��&��Nm���?Tmc�1$�ZV��#�m�g82r	*6A�q�uW��v�ωS
�@�m���Q�R42��
h��ӂS<�d^��^qد���Wbǀd�"ؾ��S�6�����x�er�d�t�b��:I�hH=5�UXήp�p�}��ɖe���������j-���|(T/���AH����5�`BS����`�}�Ϙ
��c�|ix�#�q�׮�V']�={�K7��ǡm�t�k��(c2I�Z��I���UG�P3� ���"���i�Mhp��� ��ѭc�d�L�W>�a��*i�����>�Yvĩvl���0Oƿ���ꈒ�6��c����pQ�Ta�'}ʧ9(�5X{Xj�����+Ԏ�?��6�"�QM�����`6��m��:�j0)^U�h����)��8O�_�3C5$Rby���c���bm)� ��,��'�+h��e���r�537(�.6㍶.� "E
��F6�=:���+!��Z����m���zG8ul�]]��fzOv����^�E�`��c��)����'u)��� 5�y�-	8R���X>���=e���NM�-���n�aT�#��Zz9M�Y)�3���;&CȥU�r<�,��< h�,݅
���qG��[.uHm�p�U?v��G̓��`�@�E�̂c��Ƀp���VK9I� ���[�+Y�B�� c�����U��XEvl���}�l��^�k%��h�k���AJ���gĶ������.�e����mĀb	��Ի�%o}�@��K~ ��1�P-�+����eA�������pLY�߲�޿��K��$��-��-E"��c�De'���޴F�Z{����ڸ��lBE����s��27�B�P�؝P'�:%�����c�S��j�ȡ�K�fk�o�K�\�)���4��W���٬j'{�5���ע��ۻR��:bh�ӕ��م&x�!y�{#��JY~S��O� ���ӡ�p���O��^ȗ��œZ`��%��o}�~�L�%��tƳ4���w��]:um̧DYP��$��O(ȝ�/�|����?ڰHNC>:�M�rB^�8h�VB�m�GMC�"��m lx�nŊ����"��@�_t��޺pZ>YNx���lNg^��#��`��8�R0�E{�\�����,T�����ʭt�ޔ�a�5L{�k8�{ Ow����qy�\�-Rd�@d��4ܽ&�W���+���:>~�
�4d �͔b߄L�Dz7��U/v|�f���Y���i��NA��>�fM��i*�9�N�������t�d�=�����c��o�3᝛y��cD<��3�	"����k,�������G\��m-4؎^��6�������}�zu�0�I4T)���@��
��A"{�[na��;ه@�{�y��_X\1��h�WuP����ʥ��A�YB�B���w5�����Cos��'�wPb������R=�Iol"_k�5�W�:x$
�w񩩗oҐs���*����=	h�8ʜ�-���+3��n�_*�����6_gN�����W5<�e�]c�Q��(�"v	�V��w�:h���VJu1��h�i,����PJ�/2����<�7���=�"?���{��(�����V��9����Z�r��H�b:@��uTG������H��{�����"3
�le/�Ok/[�KO��bpic�R���y\z���w��l ��%�/���<�q	%C��W�S<R�c%�s�"�j��&���vk�.M�^��Hn�����U�R�<���>���=��M�n��l�8/��X�ޅ��,E&��@q�`����~XU�2���u��j�Y��b���
�F���I�SQ�2[k�JX7'0k4`:gN��ޒ�|?E�V To"v�5˳5�7״��k3���&/a�Y-�M�D
1S��C�8+�Հ߸��T�v8b~J�Vi0��^�@�kҵ}�:~Z����fn�=.X.c&v��`I^�Fq�se��;��	�N?�65^^o*|hi�p�Š%'��:ж����I�"��T�+[xh��Q���]�
���\De�v[��,j��(D�Eʼ�ȶVXW3�L*e��){դ�n+d� �/�R�U*yܼ�Y4��d�z���&�,9��w�v}��V�?0�:2��y�XWҥX#�s��F�d��V��`WU���ٌ����&lHߛ�'5�ʋ���	R���ҼͶ��ɔ&�޼0� :�pu���������ЍР�C����梸L*T&u���S�O�t쁯����^b&{��B��|�y������g�ڹ>� ��5ۅ��8�]餤SL�?(Me{�v�t�NJ>>>B�?xF��#\���+��ܗ���'�;}KUwT��/��?!�|
D��=��yFP�Nx�<`d/���=J��<@���6�736ݬ�K��]�G �!�>��3�{ᡅ�K����]�mb�j��S:�x	���>�M�dx~���'�d�޺���K���f��0�SMav#r�:���sݷ����V���Gb����"��6���ԗ}a) ݕ8�GQ�m����y�&˾���K~��I�]��M\zOY�.;�����?��Ge?KBRp|Z���"Ԩ�t�M�x 8h7�Ljm�h���1�7(�Zw�{3�݌�Ȝ�8K���:� R��u1 V��5�U�(�,R�Q����k��{����U"��&o㡄��"�h�%a�)���j�-�J@�ev���wEC�{����9̊D�ϣ�]	b�e���\1*�	��Hd6��2 �w�\vL�T�"���h�W��}T�=Vؒd8w�X��ا���y����M�h�0��IP.H]1i�������1�&g}��_�[[!S��*4��J��m=���� ���	�G���;�{L����O2���HJ��췁M�}c�z��N?�<P/LEe ddbփ���n�_^-c�8ܵ�,�z����QA��)Ұ�푘�J��+ J�4������R۶{�B�z�C��؛�I(�V3�\�셌j�S��+��J�+����%�ވx׮˚���?>@�*B��29p�wݐH�K�-Qk1�RϤLDː�r�����L�"�Ӎ/y[���3��}�ET{�{�8���}(8������M�+W�C��.mF�/ݐU��ـ�3S�_m1���\uK�
�fG�PŁK�/���S�y��Y?/:ۨ�ѫ��g���D�$����{)0�~l>K�+-Bf�Q��֖�,�)�z�R��S��_"���Xжr�@��l��8���=����~X����߽�T�/���Ge�
���kN�=�Ss.`�������6<}?X��QY��48�����n���C��w�F����`�K�w+5~�Z~~�����H��E5%ǈ܌J��=��'�&�����`��!w���t�A+Q�t�l�xz&���`;[��x?`c�hBf�_�e�K&S9/.�*T���r�f�����w
㊇�������u�dy��T���3aq���l��@�~>N�}�v�
H�H�W�p<m	>p��'���DT�G��cY��\؂�Ž?Xc�@��u�,.���l����H�b��k����'��I1����%�)
hM�O��nɪ�x�a�OD'+XQ?u��l�^cHv�|f���ƿ-e;Y�^Ʒ���Y����h��#�&�sԭ��_�Yl&f`�P�]]��Z�Qtd��f�IR�n�C����Nq��Lɼ�p�yBaW*� ���\�( X�?q��'��O�_�!��)�G ߇-���F2[ �/�������r�%!��Hy���������L���.���	��m�kF���c�跱d
����:8-��=��h�A|~���d��S��D���<n)2-
�PLu�%��J���e���\G��&���(i��M���Q��.@�W�XZ�D���Ò
��P�ş����=�l����d���c��6Z$ýA�����ё������b�rn]ud����r�/�?��(!�0��}."8�j�O' ���ph׿�TmK���Z؛:�>]҆�χϨ$��R
�$�r.�r�!���u/!;�vt�	N6� S��\:���%�A  ��,t�N@��i��32e�1�o΂O�NX����N��&%�����-M�Z^��WGmg�	���-�L<�k�:�Iޙ?��iZŬ���J�:�(\�7�Fpv�}v--�}X��<�� �u��4Hj!^^o�[��'��_���k{<���C�?mЏQ��Ŋt;��~�Si��np�ˆ�+�33����W��L_wŗ����?���F���ףF�%�)-���G ���@�T6fC9c]8���`hԎ��Q�FH�y�6�g���*��u՟'"L|N���4�_$K��K�����^R��>�/0x������!�,5������{)�bH}|�á�B�R5t�R�G��G%q��X&�5��i�Z��p
:�(�!֖b�`.��=$*�<0ԏ�P��bL��bKΛF�2\5�al}��t��r���*����e?B\�b���1��۾	�Ko+�;��$�ZJA!�(�������|�؁D�����c5�w<��D�Ư�Ft�`F�Ϙ�Q��BTw�N�5�ݷ���K n|6�N�e�|b|�YM�����^jY��Ve���5�j���c0�j��B�a�f�(�F�R�#׸��i�n���^X^��~<�"?d�������`����%�pV&(���֨Jnc��Rdt\�X"7Fa���9��M�P�k����X�:n��v��7V+��i�=ߔ�N���W=�7�Ո��N}�^��4�a�2!�gOP�,k�.��8};]A�X��5����<�\���q��	�����;KJ�W�j0^��ޡ�JŎ+�`��1f�1�pK!�$�9q��sm���W�[�?Q�EmX��	s{`T�r_!9�����R��,o��h�$��S�s_�o��J��'�@4�c;��&��{�`�S�v��I�{@�5�J2 Ij=�&�=�HR��4�Yq �#Y-��������å��h�6���Ko�X�EFŮOpz���~-^���D
��XH�1E8����=�\���gt�L?X!�����=~��5!7/�	&��d\bMy�y�Z>�х+I<ԇ׍{*V�O,^�O�.砲�\r��اN�F��9�5f9L�RH#c3��|��5��xȭ��(��A[�p3N5IiW���K/�����
x(��>��f�肜�����CTx߁�s�y�A(���"tՇ�$�1楯&R��{'攔K���P́����#i���*D�X<�R@�8@mM�:�D���-�zZg�#z�q��wF8���hW�gR� ���~��.�Џ���k*��kW�����c*���-���Z�Z�3eN��\��5�&5��Pd�v����ozR�����ƊɎ�K0^���G��#d�z���ȠWI��-��wp�F����W��A	ͷ�K�w��z	Y�6����?{7��c�ɻ��u����-kl����3����:�\���p��rf����z� �|��Q�VN�fC��Y��}O��]�kW]�=e����6$��r�h�T�&�j��@� j�FˁB�D ����-�����]�������4}\xYԻՓ&��=�\��܂��?�$��CX�ť�P[�o����Y�Y]�*��1MOW<fY` UY���mƠ�J�G
g��.��q+E�L:��"��=�zS'=���* \�K�{\
�Ur��X��Ig1|^�X���������8�A�
���_W>��;����{��>w!c�\H�^�������O��Ox���T��y�BB��?wA,��$$�&��ō[D��Qb8��SK�k������F0<�ЌP��ݭTV���t�WT��iG }��3Bo���a����)��=1}:�b���?���zzW>�=Z2;�*���d���cU��׃�y��T��ni|���bx�� jU�ۙ�|�疖>�^��|e��~�9�,T��MBk:�w8���T� 򕖸.u	I�N��9�Ȍ��_O��v��(1ė��<�i/���<���	��C�o[� ���f����5/-}hB���P����o�5,�LꢔT<��r�!�[�Z��6%���ꢱy���˨E�m�S6_|��v�
�4�4j�R qvK\
�w۸�2Zd|5�lx�P��/����d�3͐��=}���.���n�iͣ��U1УX]��hgz�v��7Oe�M�>�"�iS��l�_$�$��	��	JS�%�����g�0��"�����e}��DS�ٍ�v�xw��{�w�� � ������*�ܘ٘e��0��6w'�m�"���8��4KC�Z�	��vf�(��qm���Е�M�[��jC�^g7FaU�Km����PEM�j�c;,�c��f3�VR#Z��PuBT!ߤ���řM�J_�h�Q��sAQp�MIa/�o���n�~6gd��Yb�(��)b֌yb���� �����yao�����r�|t�W�E��#Lɥ�N�֩)]U����c(��XL&�?��꼩Z�s镕�X�Ӑ�V^Җ�
�U�L��k����3��2���uL���b5���G�rH"yH��MYePs3��><�a����10�iF��J�g_ ��ݶֶ1�'��f�R��2t���p��x���w�znb?q����o#hdH����F-\��v��� �£e���IӨV ����An����F�W%C 0��5���R PP�8/1��{S�`m���]����E��%��c�L�/�Ao ���#nD8� ��L�T5�	�k���J|���Q.~��H�&F"�?ͥ#dB��X=�Y�̍}d����`�m��*X֤Z~�Ô���W�E�g�6����9�y����dY7�[�G[v�M� n��f��>+\�x��3K���QAd�_��n��b�' Hv�Ӹ�kԷ�F��I�H��W&����B�c!��%�C�CyŒz��Ղ-�~}ӝ�۫��C��lA�ى+��j\Mi�&Fj�?��b�a5>���א�v.O��@C�,�g�yZ���Ĩ7F�\{p�q��tB�vC�I6�^�����K3\�f/�D�>�"lL��M�G��h7��C'�d�?ACv��0�kqt�
a�h�9wk�踢|w�XN��&�_nQ#�9�%=�l�m��ǀ�0����w*J�\)�k\��"C���T�*�`����}�P�L�H�2 ��_2;E&pv�[�/���U.�A'���2��g����:5�JX4�`�j�7�~qWcڐ�Q#�r�XJE輘��s{VO�t��������6�6�9%~��2Pؖ��Fe~s٠f�v�����k��#9亣K��+��L{��B�Q>e�h7�G�CaI�A���y���}K��T(���M�����H�m�4>"պJ����[P���]�m �E��7P�kL�(A����TU�I O%*�ˤN@�#i_�ތ���$5|��Խ�K>�w�4lχ$O�+/``����L#�-�AA���RU}��y�>� TAb��0$�M�`��K�A�0��
��pZ������"���Np�|�x�X��F���q�b�M%	�I�E��EX6Uv�,�C/5�@�G�����U�2
� ��(ӅuoPn�E���呡4�P��~o
t�r���Lf5@5&����M���T���N���<���aP�]���Zu��X�Ȟb����Z#O[�r�vα�<��Kğ�?�z��{N(�H5�b%���.���_�)K�ޜ��FH�sy����a�|��������C䍫3�*��5P�hy{!� WJG�ezS�>23���a`�=5�,"��t�5��(o��`�j>7bR�K=���Ӊ�FtC
o��c��.ըy9��]?�y0AC�fH�
lNs��o��Ǐ��4�.��w��mW��̳B�<${�s�$�'�h����|/��j�����������=8�^3	0$���\8"�T� |�^��⿗&:VJ�wd����~3M;�"I.�J|>�dN=�mgaA@~36Z�˝��.xR�%S@�w�B��=��&����&�2^��I��M�A�K���l�� ����ѸQ�����m���S<_ &��[�mȍ��?�[�ٰ�N�	��2�E�*�����4��g�G�@�B��VGG�R
0i��8�=�)�z$��
U��K�8_*,�`po8q]L��e��6{��+���Q�'+����r�"��F[}C����0����Y����+}
?-[<j6���Rj#$�/s���8�0��X���aGc����zg9IY��X0RJ��<Xn#���7,48
��}NI6�4.gL��j�2O��@.���23��5��(D�K¥J�	��B8=�ޫ��k!jA��cq������s��%�4�Z�! GO��"����+�1Q����Jz�F�:��_�$�������*��X��@��jN�2P*���.��"��`r���r�'��_�yEq>��t��.�E�PϮ���r�*v���X
%cG cut�#ҟ}
S$
���v�K��IAaEd,Z��sN��E{�k��n7]�q�NH�p���}�C:��aM̻f�o�'�z���ӧ�XھUY�p/y	P�Z�̖�9&�+�c�I�*9��0�؄3���
���:q`���ߧ�A_����Ѿ��7P��]��^�r��|�5s��}znW88�\T�O��#r)�����Vދ݄YyK���j$�i:�\`��a�^�K������Z7{3m�-$a�E�y˖ʹ����P��n��kҠ��%Tߋq��5L-/u�.��.�%�
��"���R�Z�*��� SC+�}�"0���bB��Qb��O���;���3'�d�e���7�EĿ�;
�5�?��8+�}R
���w���|@/���|ః�.7E?e��v��o�,셛�L����{h%���L�Y	Ir+g�uy�ԺV౻Wݎp�qG���o�\X�lQ|~xj�"�bM�\B<�Z�[c�
h�����^]BRb��8�T��N�e�]y冖�هs��Y�"~hn��96��{/y����z�--�q�
5T���oP��������7���N����=��].�T@S�:93\��NB��KJ��^L��b�Ҥ�	)b̪$&G�늻O����C��r���`��0���X�^��Iud��� \B��t�#u��l����˯0"�Ul���Y�_�c�5���yI�#>�-��4D�^,��1-�?!ρq�М:Eޓ�A)�ݎ������^Xp���ku�R�>E��׾/Aڤ?�Q��K����=��d �e�����ru�g���PN�L
��_:���ݼ�o5'�8-��`��zZi��\�@����k��ҟ�%_���`��=�/$ms�P"�ch��v)JYĦX5O�p���
3�tfI�ѽ{�LJ��\H!�Ec#�[���E�?_Z�%u`�2z�n�����_�w��Z���N;�6��Q!
�X��^���f��U+ÜǴ��ِ/#ˌ!5U�vx ��.R��gqYY�G��U|�Q��㣳���v����������E(�R�уJW&P ���a�jtE+����D��6%�S> ����7�\�v"o8���%��	qCZ�N��l���-AԶ��K�>+p�+��A�jY�K{����CFX�Ѫ. 7�?���K������Bc��q~mU�K��^�v��'� ���4�S�Vi��o8$'�/���WP�'�,�u#�V�#(�f6�b��Vx��?���2Bn!�0F��7�:T���ފ��ve��i�1�W儤�1�T�R��}�Z<v���7��b~�*�G��я����tG�LB��r�z���Zr4h��؄�C%cb��4�:�	��;
?a��
ǔ<�0�]�.����e��{����,x�U�M@1t��EZ�p�,�}f��t|_�@��*J|QPP��8�\�㐿�EyBRₘ�%��v�ռ�?��f�2�n����tA�J��%o+����č_PW��sΧ}Y��Gz"���<�.������<qc��%zc��e3��3�Pf.�3J�w,S�S}2�' Ь��v2�ݹV��=xw̼d!�ړ���0k$Mp��N��ݠ��J��종M�������ഇM�ȓ�c�؈5V��ͫ<��U�'D�,"�|q�ng�E%���	��L"���ɤCd9[�����xx2����x��V��zђ�3Dk�dû��`�1=6%?2HG�h���i�gG0����_ĩ2G�LxV=/�)�s9��Aڙ��P ���DH?�/&�՜�Mh�/q2�g�W���ĸ�<��s���H�*�;Tn���G�Uh'O8
���i0d�<�d�dUG��º���2�����-w�CNL�O�ř��5�m�����:w_0/+nu���AA��c6$���\��d�8�@*��a����Ӱ>�d�Ϣ(GÚ���i��#�y�`5����_l���yR7$YTN�oPb�F�t�\:�wUQ�'���7���]j-��.�Ԣ���<����O�,�\�བ,/H[s�B��Y!3�?B����ƻz��G� YA��_��]y�r.rc�#^	��g��]h�L� }ٓ?�������9�y�W����cB�j{*�PX�H�0U`���V��*����b�����dZq��/��6x.�q:���F׾ル�ߋ$����,r�Ȕk��J���đ��^��k���3E��/*��Մm�{���oxLDbJ��*�Ք/Jc�s��&%�L�(X�n�Ѡ�/.��Fs>z���!"jE�=���C��ʯ���A�2Zq!r��1�2o���r2@ �-����@�-��1�yi�dk�XpKQ�F4��k���t�������D��E	��a�F�IGʽp2��W�xγ6�%��7�YƉ7�b|�:�Jú�,&X߳&�ϐ�:�ae�.�W3ƴ����{g�^,��b��P fr5��o�Wfs�)��a�
��c:>̰HX�Xzÿ�P�0�� ��j���̰9u��=������6�[���ß>@�Jb)� 1�ț�|����Uf�+�$$5e���A�S�r��r��КJ�W��ʁ:����w�oh�NF1)�N�W��g9��3(�)�fB�FE���_��F;��*�Oc�X���̤����Do��]$�R��)�
T�|��k�b�<:��6ł[�8�_�����a�[����6V��K%o�Tֈ	�M�rH��-����B��:�k�E��g
]�8�5dC������Ҽ��W	j����-h��(��֐�#Ts���#?n2^��~��۪y�/ӳ���z�9"���H�\v5L�3�e�UiF*�gcIb��nV�.��]��J �V=�i��3Y��� ﯛ��x����~�	վ8��Kq�E�r3wЯ�F2=�B�5u���	n����=��<�c�%�� ���X�)	��/o���(̪4�� C(mN`�<��&͐2t��?U�5)�띋� �W�4N��%O�6������x����0N��N�G�L�y����Zń�>�.h�4]R��p���D������`~��T!`灇JP��U�o�#A����"�!UX�gy��5�x��a�MZ:�}ގn]�:��`Tɯ]��q���ф��o��F����,��`�9�;[������i-�T`��ؔ������T<������m9GPK*?�+ˁ�	����H��K��M�	b��F��oɣ��L�b���
���0!̴>�X�5)��{P�A���#49*�
B�U��������w�zyJ(�̷�*�k�<�)�2	�q��B>���'s��Ͻ��*]��G}S���MtK��#C�i�S���Za�*��D��z���I?ە)_o����Ϳ�ISHH'[%�6L�t^��v�5�8Y��$r�n�V݇cػ�S���cu�<D���p��n½˘r5�l�۰Ѭ`�)���FX�$	M�8�WP�/f�l�T�.5$X|�g�O������He�۱�~I?s�'�Y�]n�)z��z�3�:t"�u�F����@�����(��G`(4o�9G��Ƴ���OQ��Z�vMo:	�\yC�)�������3�y�XM��>w����v0�J�g���Z�u�P������%�a\��0�{]g�#>��+�[S�>}R6��<D&���ӱRn (;�U��|����ڛ�R�7�*2ݱ]�88���t�=DI.Z������2 �T���dUp��W$}�ϚV��Y��0B���ʧs�#:�i�a>�=�i�&a���5�Z����t+�l����Я�����눠#yC�x����Ia��WT�Ǖ,ۃ�Y֢�p�	�l?g�C:�kϲq�Ur���l�5����G�\&�
{
=�����H!�h�0�~���3[i�D0v�"�N@�`[����f��7��
l۳��x�B�M&Ɏ�l�0��f�	���\�E��
��~D����cre3᰺Y�I���)�[��B�M��o���71��w�Y�u�/MÛ��P�����n���/#
�ӣ(�;"V�[���c�D�[�D�Z��~�P�K�59�{t����A���z	�hL=f��X��5E~��L�3����6�=� ��Y�Η!i<�R�4ߣ�ݶ�Sc����7�[��|�t��-���E��0�0sl�Ƴ�����"{GqݖL�Q&���]v��y�w��l��Lp�t��̹�a�m�Z��S�����������+\Z�b��ܚ��a���P��
���.�"�x���tM�Q��5M����-6��,ei��ƾ�=�\=eǯig|�U0�4ڂ
ظ��U���k�>�z%�gQ����t�2���kR��"E]��� ��A��ٱ)V�[�V2�y̓]�����G{n���r"jBWYH�p��0�eS{Qb��,�*��������J7��:�C�>���X�X��k߃�C�T��T��C-8W��h͇N�}� o�l�^a��N���|��N6�����՝�\�kX�����'H��Ҧ|������T�.m����������m��d�K�f���v��]	i�D_��)g��P^�"���:��K`��v���w���2�݇�t�ʲ���W�7����?|O�RE����7+#X���
���4b3UY��E�T_�mm���f����+��/	�ݣe�R�V�"�ܐ�Q��BRZVE^��xdZCKץQ��L�yK���CF���&��
O7 >�z]"�T+g�ڒ�Ys���#��!i�HK������ C<6^g��5�9����?��ך�L 6s�^�;�-����-��O=�a�sYh����� C~h"��Zp��WEsK`b�E�����э\v6�q8�m ���4���4�&�n>�vo**�|8U���;�-��ۃ���B|���96�5Y���׺�}�I	��#���a�4�9^��9.�{^_�lxT
Z7	��ɝ�C�W��!�!�5:ŏ0��I�B�J��8/��$]dCb�OZuf�n��#F��s��N}���d�b1<�rg�8_�43`��5�Hf��v�R�}�e�&�-�������3�,�X�dM+O���&��*�S�����E"V:���֩�Va����H�z62��y-���(<����F>@��(����֡��,%�J��{e������@�巼����G���v����k�f�'�x�*��Ģ�c�ď�z䥗C��%�W'��):�aX-��ɇD�;l����U�	*��W�����}|/��5$��5�/
�x<����A���/a���O����3j�Ⱦ�"4�3�7�������D)�>��|�����+�Qd,�۝�>���������'-HM�ۖީx�<�"��uκ� �A}�)N\�M��S�]+�P���j^k(�:�z��)�����ɂ+<�]�o�p6��a�sǳ�n�x!4�pp<&���OYٝU�I�a����q�f��VZ�I�Q:��Ұ>�L�*��Ac��sA�]q��-��q�m� ��5��I(M�s�8��~׸z��7��wo9/�I�?��I!��W��n���eUpZc���]�a��ʩ8D���߾�jh^�ֶj�@������w��r~��3�B�{%=5x>���V�n����@����%�)q�'��7���uԔ�)�B8��֔!V����m+�{�m����x�h;�=��=�v��tY��/��6Ȫ� &Wx@��)�Hj5ϣ��j�i�wk;�&��`�������� u������d9)�-:_����=B�9 saŢ�ec�,��>�h0�tf�����C��s5�e��	g:�i�Q�XW��$�M#%��؛N���C ��U �W�J�-�b�W���-m��o���/z�5�T|:k3�J�����nkހ�X�EڗPM�=�XRG �쪹B�����'l�-	١����*�f��RܜuÞq��7��c�4�?��jI�[/H��D>�5?�g�x�RIs1�W������g�k�a��#�B�s\��"�������E��l�$s{�u�ň���S��9C.��N?��}�oBC����%�B�o���Z¨��ڊ�֮E�,�s�	���M��	�	�L�Cݑ���'ZA,�8��5E�P����Mॊ�݀�n٭�損\~���0���Z[�����=�{����J�}��|����-�������}ETM� �#!ꋥS��}���`(Tb7���
u���$�c��_ld�gVX�jI�L����*i�ӯ��Q?0�Td���m���*��Q���Ͳ�T������m��?$�+�7��p��+ͷ��Ӥ������!��e���;�i~�3����ˁuͤ�$>�d�c��_���@��~Z���Q�QS=��.c�-�LФ�ti��`��>�E�{��}���2��2�16
q<[@�2N��/Z{P��`��ax�O�i���1�T��R7I���%cQ@濿�s�{�3ܿ*J*!���X�����S��(>��$����`� ��_�LY�M5��Z��b4�"�
[h5�8���)�l�b�!�qS�Ԓ:G����Չ��SDԼg��j��/�T���ov������H5�<�?0j;��6�c=�Aϕ]E�ܿ��_�&0�h(���Z�ݵhu"w��}w��1�F�ȭ�2�ծ�SɌcj��L�3�62X�T�~ci+S��nB��N���?X���Jƕ�O~��u�Z3�-v����6"����v��Y�P�}���&�tn4�~�oݣ?����L1���f*��s��O՛�)����0�qt�g��Ռ))��L_\T�`�]�e��`_
)i�0�j�md������֥�	E�з�B\S/U���� �J���h��0��a��қۋa�ԅw�i����~4q�@=l�1�%���/�tӀn���g�j邖��+1ׅ9��r;�:����_x��w�]�_Y+�����r��}�fIW܉7獑R�E�ŅMq��q�*�nuw0� �]~}���d�hG��^�)����75I�";����@3�H���Š��k����If�P��˴?*�9\���r��^b_P�T�>0	%��p��P�h,�j֠ȯQ���}��h���W�y$��1鏏|C���N���pn� J�^<8`�/���W��:���4�.��Y�ka�{.��a�R M�D�y�Q���
��oh+L9f9F%����ޅg}�^i=^��ݎoƜ��f=v�5G���_���}�'���q����pJs�ݞ	�Dz���[�����6W���!������.׹[�D��#���ֺ���*"Pvb�.%H�I��fo6�(<�h�u�MN_
g��s5!D�V��r���8�S�iʵ%�l�$z�����G��_�}�ȸ��a�ddu��z\����vE/�(�έ �a�Z{�_�}����%�jH+2��J�8�S/��v�"P�I���K����S�h�;S�sH7q��Ft:!W���z�I�B �Oh�0c���M�"	�
։v�Eh��l_�+Y��Y��Ǟ�,�EI���J|��i� m�t�»0��<��/��[����B�+�[mEg
�+�m���|W^��������h��m�'���v�O%X�K�mQ����>q,k�Q_2�_�E�<�C{-O21#�5���H�� )�ַ�`IF'f�X�^>	XJ��.8k_�4�~�1^i"K�(6hZ~GT��o�`  Ƈ��6nd�W��S��U<����L�mȬ���g�x\P_��j"�B�l�����.�����|U��z�u�UnD`���9���aa�N{�a��!�ҋmXCf`A���/a��+��e�y��¨4�X�@:�^��Z�DE5���f※�*5�(4Ж�	8�Y(^�j�C(��҄�����j�gK�Y����v�^H^Q��!��t��UA�A��h�B���C�8�k�64���aQѝ�@1z��sI�5�N��|���	��>b��owMǹku���X�A1u�����.QO,���hu#��А3/�1�g��IF=��X)�y0�נ�5:�v4N����bs	vX���!��Y��%�bB�����$<��2�)K.b�VM������[c��8��^��8��h�r���~>h�0FH���P��v���|gj~�(�(�V"n6�
:��:�>�Q4��]]U�"��Q�7�-�G�������ի�~pPO4��{���+��@�F�D�!�<Pqk�����;� ��t��-cG�n�+$��<ӡ��v,0�e!��Qn@�a������ޝ� � n2m�2�� �B'�븎n*@�@Fb:�>�P5W:I��A�����Y�%�4�bK�vU��R�&�b��-3�;PK�̚���G����r�������g�<1��U֌���|Ge?-/-^IbFC��I�b �wy:^�*�Y����,��(��ϭ�M�2\J-�s4�O�����T�T�kL��r�M�����q��;Q�<%���m�	m$�M��
G�5x�X�K�Ҝ��7Ӫ�?|@/_r�"�KDǋ�F(�1���΄�K�C������ƃ�0?��V�ڨa��1�W7��K`��$X{S����T�	�k�$" R��E-���u���{�:̱
�~�O0�}��h[�W=P��R�E�A���"i��̴��]��vDJ.�j#J�0`pВ�luL��X�ϧ�x3=q�d3�L$��;0q��U�7�y`�>���I�����H�(�X+��,�����Ԏ�TK��?PQf�}�W�pR?͋s�6KS*6BǤ�}���. �V<���w�y�ד=a���_@I��7�ԍ��9+��HkW �@�H;.Y�T��ɯ�dP��b�ܞ�yP y{�p�ްJ��8�6ڭ�=4�#�Ŋ0�7�̯L�Ы��i��*N�i�a}U����*�R���SdXݍ�<�)��cW���P8�8^L4-%Z�">����\�?)v�:m��6��F���1��?R��9�=�%����
"Eq�#��ڦҷT1M3��I��!�f3J�7h�n"Ɯ~S���@��f�S���y<D4|iF~�
t�Qc�G����}y���̢#y:�V���7��`_,���=�kY_�6��3�k�s�:���J��e`4�?L1��+{��B��Zb�T{0��'��,'�r�2���r����ˈ�>sF٥��QT�>�ܫ-#��P8B?dᯩ�(�ҹ-�(����d��]?Մ� 	3F	�����[/y�D��a���w:���͉�n\�A�|���?
mh����6�=�Y�E�8?uֽ��*ʢPc&1�����Ʉɰ���q�IyTK�dK��׷0An����p���Q��u#��SF�
�Z��L%Y��V����CKYMMV����|�)���,��(��+�x\՞@��Ni�]*�?e�CN^����)��ڧ|��8�r^��	Ny�m�"D�8�_�9��Rwcd �J@�3��� R��=�w�3��j�!S�G�n���,��������Tp:�8c �_r0%l��X8y>ǛGm	�v�D�D�)�vP���(�#�}%��?ϱJ��t��Z.�����R�'�f�yɞ��"C���<�f8/����(�����W+sw�{N-<�s�Ў����`����i�񡯨m���!�+c�`�2g%�~R�ڴM��.@2�Ъ4��A;�����1����[���[�+>��X�de~t ��ƿ�{{<�e��6w�-���⁓��_T�%�B�1뭫t�K��4�m�ڐ�7��Pn��U��u+8�cO����;��i:��i��ď8P_�4�E{���h-7�A�����3o��]�����C��]�1�vC�O��hh��q�L:慎�����>�������;C��f(�$�k����ۋ��7�%��` K�T9 ���b�JX�!o�C;,�K��y�Z��+|`L�S���E}��b����A�����-X���M'(��}�U�Oe��w�{fU�=+4��s��x�S����:Ү՞�=*�W��{�(Y��S$�l�t\)�gl�?*��h��BGc��z�44��op�0�[�ġ���L'��G����]ߛ	�!��B����X"4�WM�F�;׭�0���Z~K�U��Q�q�ĵ�@<K�߄�i]���K��0��B�y�&�D-s�y*���=O��1�Ot�M���=����%����i8C}���R����v�����"��T�7�He��s��bו���/T�&$@k�G���}<�>S���G�0bB�W���ե�㻓����ۓ�#���}�*a��l�6�Y�{a�O��T�y�{�s�gg�]��T�5�r���#p�{�Kl!�!HoБ~�.�{�*>��v��4��Ѭ��YF��\/)I�NC��]|<��l^mN�ۄ�_� �E�T��UʐF6�����߭�_|�Ě3�~�~#C�4�*\���Z�ϚRGGg��mz>���M#�4*��� �LB�qneD?-��2]]B��J8\����`��R�eF��V��.'3�$�S�WD�������XR7�<J�#��9����h�pV6V�E�4�f�fJ!�p�aD��Y<�`�y�{����<Ll�?�µ]�;A��
�� f��;�c�?WLQ����ݸ6e���<3_�����d�
_324�>�&l;6ߣ��������1�ZwØ"�^����*�Ԡ����@��AC:�=��Zr6��F��� -e��\���l�d�/��4/�$��m���Ke�\��,�� Rك��׏�!���<��f�|����j))��)[�q�t�Lt{C�?���s�A�6n���_�����n�s�4�H�w�}�#�W��!�RɁo����)|���yj���Ъ�1��M�:Zt�h������C��z��=�K������Sh��r�[oj���k	���E�m�@����T���x0y��U2&��w�L>��zmu�G��8�I�Z���L�34Y�ԑ"�� ��ML�3�����
�{��'��W�ra<Q���v*��
n!Z�4����}�c�Ag��n��"�M��i���K=Z6i"�ki���P�Õ���k�O��u�.��Xek`���+f&M��Y��
r9�mU�4͞�x}���:��oh�l(�"2E�nnn���1uWSE�ȸ}�&^��yn�Z{�>��9wG��ɥ�[G3tfV� ����ځ�aΖ�����	e0zMmBu	�N����&Ua~��ރ~�ѹ�C ���'�I��a�����"�C>�;z�1�Hv�j�A����5�/���#��ym�\)�3�	.��7S���ߵ�)�Ɠ����b���o�F=�!r�۱Χ�z@ڜ"��s�m�:���#'|"�溙G{��Čy� �'(j�$�'�'�O܆�����5<F�C���Ӷ��}GSi)9
 Ma	�O�ʮEș�V�
����7���\5^�GɁ���G���f��f��6"�����(Y�4Pq��7�\�`��;����i����t������Х��L`'z�-w�x��� 
|��"e$<�
Y��P���yw��^3���~eO1/N_��kLY���t��`��?P{w�҈��V<2T���ޫ��R������9�f�ȔO���V�E�6����\w���C'���
i�P��5y��<��_�e(^>�+&Ɨ���mi�S�tlV�x�ƢM^Oڵ|_�[�,-P(�����$�\# �^����
!�v�;��d4a9�|�����1����RU���a���~+�<`<@K� c�}��	��O+�'����8�w�ܩ����c���D��X�_+D��Ř!�L�b*w�>b���U� FU����8Ӹ�a9�O%j@ ��(�|-��ä�*8���2�_���/&l��9�$*N�!�u#{C��5��!E`���#��2w�&˭W�*���&������Q#U�e��`o���Uk�	����h&:��[F����)=�D9�;����ϳ�S�V�Xc�6k�`f�h�~��P��{��}a�����-?/
&��k?&�)�O�N�Pm˷��-��'r���g�.QZ��3��6�5=q�	Jj��AE�I)���*Du��:��-� �5�/RԵYۣJ+�&%�̘�~��Je���j���FJ�m���g��b =�8/B���Ѷa4ŦJe��^"�f���-�ɳw�LE��4k�x)A�d^�]�2q� ��L�H��~�c�V�JprOKe� U�E�lQ��y�ɦ���@n�Ԣ/��e��Az*Ưܮ�I�1+���"c{Gt��x�����'�KD$**j�P7=T`*��:0�z>��-߂߼�-�}5y��]@ؐ�s|�i���g���b�Vh����[��Hx��f����\��>L"���A�A�wC!��>!�a�Gb�8��lx^pA|���6lTDѷ���z�D���>P�o��U� ~�9���G�=L�g}',�4�$��{%D;l�����aTwb�'!)�2d%f��VL�f6vr\�;�*8�dl,�ߎ*�(�r���f�6T�$��˹�@8ĝw�ڎe��˹o�X5��^��Ы2aDe�U�i�����+z�)��0@�1k:e��z
k������T��K"�a�zSU�J����)j�W�X�1޻*���遵���Х��Vl�P[0xK�H�ao�b��҄Eǉ���g:�bx����,�[�KH�LL0�P�ځ���KQ��L�Ii ��f}<�9�Öt����f���'��03�O�{kd�ϡ�ц{)�{�t\�-����3�܆�{�<&}�d�H8�2�:��2��f�J-١ ��)���� I�{I�h�3�T��_fX��A�'V˨�̩��Pd��f�a�_C�p��c��v���z9S6����{j�rxg�MX�~c��f5�`����8c��/��҂���̜6<���~�6.��$y���d��I�Y��s�R��Z�<������kEg��ʨ�A	��#nv�f�4���>޽�/A��!*?t߻����^��c�h��vcn�4�;ޝ/a{'u-*��I7pvy%���������/�"�s?t~�Q̓V���r�*�,5�&�,7��Aso]Yrɬ����ZЋ�/�3�"ɬ����`�YF�\�s�����E�YL��I��g�ń#��a
�EQ�XAe��Aq3�7(v�j8���_���P]�~��B��yGk�u��Ψ��nQ0�Z.��ŁuB�'4�F�bP��M~%�(=����+u~��[�^ 1`���h"#�����HJ?0v���#��D��PF1Bm���]�23'M���?������-k /��;{�u��ڈ@�L�	�޼�^!�
� '��r���vh B��y��ʦ�ӣ��㚿A�d��L��
{�s�q��Ͼ���&f���D!�0?�"�\��߿���T��.uמ��4�h�Ea�h�<y�,������\I�����s�IM����e��mad��_��HBr:ߏ����? /.�U`�Z�ai�f�{�E�1���ɇgY�%��8�$��i'EYD�>qW[�,�.���J.���Բz����vz��h	L�Q��n+���]1��K�R�Vo�Ҥ�z� �20������˭��(4��П��^~���߲K�U-,���3љ�t��F_�z2 l�I%`��rG��{���ʅy�f.����ͳ�-�"4��b�Kj2�}�D��U7C�gH��'z.88*b/&N��x�O��Q�_��i �,F�i�� %�&3+�[0�ep3bP-~
�g�8)V����[5��@}��M��^A����`b�p�@�n.���A��� �W4`�5�jv�%��;m�E�t{����f���sz��2�`��˙���R[,��I��������O.�26�����%z�N!M9�.KO3\=:~$ɟ����>�t�kji�]�aA^F]j?��'�7���pɘ���Ug�E ��T�Ѻ*q�W�y�s����˪E���Y���9�����GW�7;'n9d16l���.�V��� +&9����iaI���o^�pף<���\I���g{9]u���U��)�LaR��! � �%���=h}���E�o`n5����=���$G�=(��cpS?)y�A�:��Jq��־m�y@V��o?E���c��/5��g���������Jb�;|�����>�ى�s%Q�SeV�BE�L��ӊ};ģE>����A�8'&�����vA�c�`�/뉎}�o�7��Q�\ZD��dy��M��T�M��_�?���~��,�����
w�AJ[*x41�����!8C�T)���V
��ya)!|�hkXV�#s]�`XW���Ds]QR��8�w����#W*0>{�Q��W_�"#s����wv�` ���-�� 's���9�fZ5 G/�%�`���<`ݷ��R=�Q�+��Ph-���fA��*3���@�?wk����3�����V��<S�:6m�ձ��z�7 ٛLp�c�IJ�@��C5��j�Ѥ����J��_��t|����X�Ol�4��c���[��rH�v`ж���,ӽ��OP}c�$m3����R*�Y>m%�BSZ-��cƪ��`wr��X>��0�`����ȴ���VZM��-�?������ji������������#��i���/bB`����h<Oo�!��e[F	<�������һ�f4!؀H7�Q���A V��N[��@��o�_��lVd�а�ͱ��'��Q��D�(b�<�S�*ڴ�~���	텩G��Y�{Ub��{`2��B6&�÷���쥻�\_�_h������-��s��r�
�
0��]b�7�j�ؽ��eV �h�6�������É�H�q�~� �c,A�̃Q�i���XgĢq�����uX��_���:	�:t���&(��[�E�ƍ���v���^H,�O[�}��-�0Sqh��Ob�FF�04����5����B
6���#7�����,�%�C�k�c5�F��b;	`N�;L��ʎN9��E���ҕ�]Oު�M���]@������sW1#�<����+noi����L�&!Շ��i����U*�B�`���Sh-c(.3j�(�+��V��E�S/yBTmׯ#�q���tj���R�U�/�j��Q�:�w���;nIm.�|�FC�&_61H\5��:Sr��tv V���ՐѯC��"�a�	Z�ep�)�� f2�^�Q�(���>u
x]�Ox�J���	����0�V��!�����6Ij������~E�@��1��*�[dճƥ1��x�R"���,�����Z�h�������e�ْyYq��2��VB��0�$R��-�Osc�R�w��|g�:��vd\��JB�����Dc�	@����W�4�� 9�O9_���R���YR0Q��{���r�T旐�9#a�j.&�zUХ�}�8+/Ə>��"��Y��~�홖)���Ў^7�jc_�������R�?�N���)s���g�EZP���%���&�H� ����S�@���[9O�v&
zt��@��C���5���vKyHq��E�>��%�%�$� ����0�)0O�(��XK`��ü-��������F�WX�g�W�v��~�(O�VG�*�\ݬ��m.�q�'��I�\�~eKM�_��:Ǵu��[=��5���gb�O9L�ީ������� �Pw���V0�i��_�X�Lз�'듁c�>��d�i����cb�����v�ɍk���-��wH�d���q;ɒ���Ȋ���r����5��DXr�"PQV ຤�5 c7����z�C��#�(����O�ý��QS�gA�YW��~[:,&�f�1')L��`i�7Cp�T����X�+K���L-;��M�6�w^���ۃ���$�����UD����?��ט�Ve*	˷���Ru���ʾ%� ��o	�JUa:IY�W�T͆�6�埖��N�u|n��XZ1�9�V�m_���ס����u�s�=Z��.�����g[�Z�kI�蒤��魔	n�9���RJ~Ν�c~P�"����lE��'dﮕw5���M�n�i
���Z_@��.��+4+����=c����NYf�7pQ)*f��y�O��s!5��U9�ec��E�2�6��a���\a[�d}�����)OA����[g���(���^���y����7cSA�z�BK���p�������{�M�dRv��tP�О�/������������������pj�_ߞ'��2�^��h⚷]^p����8�mW��m\518S���EN��Y=_U,*��B��͝��Ő�����U����~s��XSËQ�+6��`��������P���ߦ.%[��E�ֿ
Ŵ��#C�(3?��j����@�'[(�L���Hmt�P$
�)�e3�c`��͂��
j]�T�~62cy��eS��������*�[���RJ�;>�n���mjŵ�7�Z��{YgN;�-�������헰]��ϙ��@�!�G! Z:�=C�]����!����K?�e�:r�ʿ<d�0̨rr�����,WdPk)�XR֝�q#��ݜDe��lד��r]�}�FѦ��(
y,F�%d"��m �vV�����_I?"%Ip��$"2���^�Vu�=&��Q!� -��D���M^E����I��"O��Ct�٢�_�.�%��3m�����c�SKOK�7���ј�,&�+j��׶��Է������� �B�	a���Wۧ%�0�Kw_3�yw��)�>�V�W�Og��q�E�� �,�MS1e�""S����M�da�=*�BXiF�|ӧ�fW�$�`�<�5��J�P�W��ɰR���5am���P
jDi����_Mo�\�0X�!%!����'py^���㾠��?�����7���ԶRf�YƁ�Z0�ғ��Ў��	�K*�IK+w;�Jp�XA��������^����5��'��g��'΅��G��w���ey[�K�h~y-E��|ɽ!��Xowv�Q�`��>��!0{f��7�戌�r7 WJj��v7��(�qu��J C����V��&������X�\l�	�e{�\Z�2sÅ������1�wt���}19�4nI��K�t�-;z�����:���9�I�t�_��lx��d�҉�ՅL�&�mʍzӝǜ��1ުH6�y�=�{�W�ay�I ���ttD�,/���6����Ōa˱�1���$��-�m����n��`�M/����a �߳@P;����rwJ��x�(��`�����|�4	l��z��3c�5�v̚�����ٗ���
�>��>˳��0����͸9��u?Z%Y�\�3D��զy����Kw��* K;�?�@Q���ϼhP�{�!�������I���9*�d��ЁW��^EM?ʽ2�ĺ�@�J��l��$/��N�kK؜O�h`@s��V9������e���(����R[΍7�3�Q��C�IR{��,h�����ߠ+��f���d˃�Ƌ����!�0�	�C�UF�w�A�ydQ;e��N`ً��X�Ц���\���\eR�57�#k�_�Qx=p�D���R����Ɗ��E�:&�(4���&��w�M��'SEf!ę�۹���yK��MSx�m�^���w
�/D?�۠6�[��f��O�r�qB���PF;���B�Ӈ�Q$��E���-��l��7��w��3:"��\����]��%0�����D*��R��L~RV&-�I6x�oʡ}1U����>�����|(���K����{�҅�������;���-��C�����y.���)�Aŧ�@�L�hkX��wb4;=���Gq7�A�O�{�ө�Ǯ=��Iߋ�����?̴�rj���$�E/�W���T�R(��̓��@���&J-���t�t5��$�\M捜�0eR2��ir_�]mG?0L���=��Y��Cg�5u��#K��ؑ_�t��?���<48����$����78B�S\�z�*��J'�)#�i�
@=���D�U�A kj��k��;�b�RlN$6R�Db��q����-����,lk�6�?ֳ�I�L�>l�Gt��Z��Uc�jri�jx�Q%����\-����m��$!��w�R�g����lY]r����]��{�i��Lѳ>}C$���{��;��R-��w���d4�F���IIF�F5F�5U4����e�-R��}3w	_Q�A���B��3���r�V�~�o�	�~1>���ܗ'c�c)�	gF��#�؋a���!~h�j� �9��OX���P���r��G��~a��nl-�R��8���Fa��6-� �īRX���U���Iʒ�>��h�.S?����܀X�ţ#��'�&�:{=<.���-�OgI���;�*�����) P�sb��/~��^\����+�rhր�a��f��f����6�k���[�����C��>Is�����DfB�}9�e�Ǎ�� �2�i�l{�1x�i/�Uqh���h將!��#�v����b��5,b�0	�
�^�>���BI	B'������,fC��3��m�v�]�f�Y�i�p�)���|�%[�1+f1�/���l�V�َ���m���=ɷ���A����7���C��9�ҟ"Ѷ�
}�M��Y�A��l7�<��t��ul�V�x%5-7���P�`Z�H6o����c�Tn^��g�ˡ"W�C�X$y�6U\����Nr��W�i��z[R����R�jW�ߘ~���xC�_����$9���,zd�5-��J+�^P����
RZB����P�M�&`����V�ڎ�+i��[K,����us����t��2Î�/G'�xV���8�CO��M'����sdTos[BiՕ4&�=v঎�8��:ȕJ<���-h6��F���恨+����L����	�+��H�햓�>"w"�8���O.�� �Hc"�ưk����D�4K@�S�������!��?:jzHx�yoF�Z�V���9M?�\��~��}�2��?�bN]Ɛ�7эL&߁�mBM�U�O%o��M�ņvo%x{�K�[]K�*�t�[�y���WNr�RV�sK��.t���\��=</��wY��5��/F��C��4"؛7ݕ��`4����;��E�G��c3`�T�)��Ш�m�Ӯ4#�5��+�?$Y0B0�:}G�?�����9��e(1	����@��FQR�V�ܰ���+�����_u��mj�b��r_-^���]%��}�T~x�tF�ڈ_�c=������Cs|4�|���2;�0��yD�1�6���[Nh4�B�P,�	�6oc����2k���bD���`�D;ӱq
s��$��i�OwQ�:	���Q�R*�Ws�k��b�-�V�y��>�Kv��D�b��sM��D�o�7w���QDS��X�O�`1��
���@�����;���{S��z6�KP�"_Ѫ��q��ʙZi@�(5����^����LbNp��iN�Z��)�-��,*T�e���D�Kr��,�����l��Ȱ?���%��k��f�"�%G8��R5ǥ�̹��F�r�,K�b=J��-�H:�Y��^k��Ek���f�(ED�oQ��5"�~��/;\�<�}���-��D̳kD�� 8Rý9��Fz�.��͐�E=��"��|+eF���w`.��١�K�V�/��P�\,�h��u��ǐ�����[��,� '��*�>�k{ cU�L1#H�]�x���B )���fc��%��6�bi,�����LK[�J
���e?ȍy?@�.�S^�g���s�[V�V%�W��NRg��px�X��d7�T�e��;<���m����P}�ル2�ĤeH�;�z/�۩T�j��2u虙k4���f0ې��l�,a�7�G�����M
,�U��a7U6����,Y^�J����"���A�|��mP�
bkQ��#�du��\��#���T� ���IvG��C����[�;ء�>�:Q�x��:���$znn��7·���i�@���T���%>ȩi���x�}��/�ϐ�����if����FGz)bk@w7��K�utS��V�������@h�Xq[�㎯u��~	Q��ї�S��ʷ�_Uir������i	<�[���1}Y�g�x;~�d�}g�n!� (8�O	�s��=�b0��B�7��p|g�U77�63X-~������I{z6���rΣ�v�iuM�a�R�Mכ���w�E��d��O�1����4O��$����w���Ç�'��i^Ѯ��e�w�D��n1MX�7��j�(��)
o텺ٗՙ�(�w��}�x�k��;o NĄ��v��ڜ	׆Ph��Pc_�Qm Q�����0��2�����ə_��l����f#Pn����ˮ���mO�"��m�\�7�l-����P�YvE�1�!`/-T(0�6�"��=8�S��a��F��t�*��~�Ӷ؀qk�{��jmE�fY�k�bW�c ��>������p[�[& ^��?�4C�%�wG��VN��&�s��A��(C'w]���6Y��PSR@L���7]h޲f�\��>Ӫ0L�NOj}0=��1��Vt�k4���j��S�ׯ3�
H�
�5n�հmc��[k��`���S�,X6���V�#L��˙�Tg֛��'O���	�@��Dȏ��zDW�m��o�j�btZJ��#�z�]�����κ"�7߫���@���h?q8C5�	5{��t�	g�/�g�ǃ+k}�����z��%�����;6�&�#߇���&��������,�H-��V�x~L�ϛ+���nӼb�Ҍ	+��T�lͅ�;���3�~��=?��\2N�j�_�.��QI'��q���.�G���Z+�zrH�:��]�/��0\� (�*�X��(k�>�g�:���(n�|4�����|�]���	`%ݏU� �&�tnv^M��[¦�[�<��YI��q���jX�H�?F��^�����֓>�$ۈ���l�ډ�c��K)c���u�h�]8�zw���U�8�Y�YA-~�,�8S'�h~/0�|���YM[ix?y���A�?��h�5����� s�	��ޅ�0FY�}zM�4�\�ñ�M�+x`�Y��!��5;}��CM�7��e�0�e�S�O�u^�In�(�Ҙ'��d�e��������:N�S�͓�<�(z��dB��a�n9�B����C8��/�apF����Z��l�6Z�=K���yUt=�C��cG@�T������gG� �T����<-9��/�^#C����[�u�o�PuN�~��d�ޏr�VlZ҄ƥ������z���'V=mO崻�3��p�Q�d��~,(M�-�Im�z����o�7zgB@EL�t�B�i	�66@xi��� K�~�tR�q3F��_Iq[ЊP��j�����F�&��´0�� C&A�Q�p�E����*����)��o�e)��Z�t
�*��^lZuKr��Dhx�����u���ܺٱni�]��3.^�3{��9�a���w�СE}��kJͰ�����!y�MJ�=I5������H�)-z�:�[az���WSF�5[}�ךe��mE�X܆` o�"�)�a���"��dp�[�=��ij���-8�,T�cr���åE�z=Z���]G���X�fU	�me@e@Z�p2�B7w�*�k>C�k>����n��_g�HK�T���,τZ��m���#V�z���}�.N��xm�C���%,���9+O�+1��-�b�������������?�ݏ\���E��J�,�[�_o���Е̋rγ��i.;���]3�tJbQ}����,Q6��Zy��Z<��y̷���765Nh$��7�tK-�JP��cyk�q��f��~I|�P9Pj0�5����o.�MU�bﳟR��D%R�3�GSv���9p$z�(-��[;�����OԈ�=�\}03�l�����DNr�@�z�a�wN-� �M�cr0�Ft�Y��OW������s�ȱ��<�5X��g��+���8=��[�cG��:�bT���D�*E��c�G��ˏw��ϦY��.����{Ҹ�'�j�[�aF�������a�C��~�� \��]���� p)����0�[Ez�jk)�E"��#0�@1[ lP���#9��i&fͬf��P������!_����?vÙ=�Va������T2#�b%2��Io�y��"���㯎���cj���Ow˱I��{�Vv˂�j��v�_�?w��8k����/3N��M�0X0Q:S�b��Y�5}x>�*�ӝQÌ�.�*������6O�?�TE�~�I̳Z�>*�fǑC=U$<W�x��&t��j�_$��sq�x5u7j&���#*?��Rm��F|�VS��Է�6��p�u	��U�!�^��fe�� ���Go��Ĝ��d�/3�	���V���J����c� ���W���C��D3�`T_hD�Lϙ{���J�c��CR�@�~Sv΢�,�:b%��~<E���]�z��_~�o��$Ќ�lM �1�̝2w��4�}�ο悠�yk�u2���K�#S@�R��������H�C���u@�J�����m�E�����>�k04����[�\�%Ä;�s��7����$�*aS(�v���.bO��K�\�T+.���ҙ��g(JCR��k�C�\�7բ�,�PC�{�Tr ��h�ɭ���EhJ�"��*e�� ��!��f�g����O�SZ�:V�'��j�)$s��վ��������M�*'��v��Q�T�fn�O*�>�Y:*�}Y���LT��aϽ2��ա��z��e�zK�_-�&G7���y4l����U2*�5��������ĸa��P��~N�V�X������{��`��/g׶�A>N��z���ͮ]f��PN�^T��Y��[�[�qiT�{���=�"Wbf(�e-F��7�L�����t#�m^7 �H���2��>�t5%�͎'���x/�5��~����<��<{�5r�pOJa#8�Ci�<�t�8�)P���+b��\�S�}�[��	�P���Ru iQ'iND|�(rf�x����u˿ڤo����>K�P�M���?��T��	�&�z�&Qs&��Y@�Ε�k�;��nA��k��,��*�'����/2��s<!(c�K9�c��E�EAV���ƑPALߚ�I�W�
bO�%d6Jξ�,��j�����~��wM��u��0Ԍ�/W���`T�d��d��hޞ�u(�-���@�|�ʠ�1l�Pz�Fa��"�\��)}��XG�MI;�D��&�;�(-�:�EvC��]�����fgq���ͳ5���VP�� 鲇�\��K��
s B-��B��u^2�\��Hc8n�cE��ܭB��y�]d����/1��
h(��{�|B����7ا���.��Z����B���4�d�g�l��9��a��I2n1����	��pjĿ�㫂�:$��X9�	{*	�������/��+�cq��o��y�DsyOʿ~�ؕ�8�����&�#;K%�X}�7��`����&7x?��*�r%(�	�4gW	F�h�V�=���.P�{$�E�ʲ�k�Yx��8�FL�l�)�a$�͈,�b��La��8:>�NV�Yd�$�[e8"ɫ��
����2u�=d�?yŎiHԛ*�1zp����h���uI{2F1^;ň�q���[�xmp���W81"���?~BW� *&�0�UKR���ݴOU��b.�)��l����(3���XסJ����LJ>����?��҈��&{�ysڥ�i������E!��mb��O%<�
W�pm��]v}���{='Z���1��]?��2�3�}z�z�u�%���:�P_D�6��N&����b^�'��i��>�IO�\,61�6�ᓹ�Q�%C&v8�ڷ�=cd��/�{�Ml�p�g�h2 �ء���:s?��6 �a�Sp�_.Eې���UZk����b��o4e����Q���sw�)(����G��k��^���mp#������a�	Y��믫bMݎŵ�C^lNn}�Ps ys�^נ�'��_��*P�[�qu:�Rd��@7d�Cz�ɸ�$1�`���cA��܊��r7 �+r�=x��n���W�����]#d8d�Ė��p���w>����gFH1���-3z��'
hc�G�Ӯ��]V�X���_��v�w��>1g��������^:�#t�,ܒ%���F]p��x!��^f\�w޵�e!�p�8�P���*�ڔAl�ie��5��h�g�à��í�r7<%�9�~3�A�GS #$�2�v��\�f��%p#sͯđm��7�m�f�*���m0R��;��,N��8����f� !��ȑkƇRJj&�9ؿ��	uf�X?��%6{�O.(�y�����J�K}�g�k���ݵ7(&��k5ڍ�/mS�ΡJi������Xbwm���Vӆb���J�x��y�P����k֦��~Z�j���S@x�?�BԖ����9�=O0��(?[;`���@1k"�Kj�^Ze)�쓹@R�fx���S�n�`w�[��6#&��c[�\&3|�m{v���-B��Ms���_�H�|�ͩ��!��$�N}��f�Afĝ��;�����Sa��b������^��w���f�u�dk͇݇� ,%U�wįܥbE�wD���y�@e���i��h:0o�v��h~��h�T��58����eVN��h{�CM��D��N�<W��6|�΍S���E]I�nr����z�LW>�u�c�&M��~Mc������f���6�����m��h#<`�E��l�D��
l`QB�%-���%;���*Sl����l��1�!���2;wREu��f5��_Ħ�y]�"_�Ǩy��WY����!����bFAT��>e*D}���Re�������>c?�c�@��o��$vRxa��e7J��kO3�	�-Ԟ�=��֍���z|�rY��fcO��D:Wy�_�.ꎂ�(�nMd�&p����˱hn��Y��|�;�^p�?L�hQȶ
0��<��ݠ��,XҲ䩡�/����a%���S�e�'jS]�D/m��_m3�
�2�����K�7��� CdLw�O+� O���l�����"��&z����%nh�"������R}-��#c���v�prŜ�V��e�%��Q��S�L��ݮ���.������@�US�A��9r����^hp�[ �0mĳ߫]�ܥ<:APjRT$B?�:�.�D6#��t*���?K���8�R,q���l����T��j�J(E=�����C-#�@���]�PBԒ?f_U�h{����65�(/Y_��BF1�rU���ߤ����@cVQ?'{ƙ+(�� ��zD�f����A���tC �Y�\�ٿ4�	{�N1�$�:�h"�����x��.��8�ӥLE�1�e1D�n�������-6L��Yy�:���\���*T+���[��z���p6b��������S)�����IC�	V��b¬�x��^`;�	wF��F����>�.�-��w�<��ڣ�f69w;�w��
|��Y����!��W��+��ǘ�AEC�]k� V�vH����K�L�{�	,�9]�BfAG�1ᤰ�PX)�e�.\�c#�>�>��{��J6�:�n+'!�8�}�[�`��S����O�=���F2�L	��4WAV��Y�R��ٳ��<��&>��l'����9�ǽ>MP�}�R�]�"��ASgdG���g�ļ�oo������8���C�݂u�WsH����͈";�ȡ6�7�rC-������88a}&��<�B\Fob��Y�i�]���dޚ.�f�f���������.��Ѥ�%����C�6Sj

V�` �iR&��f�����^;���|���GI=>Gt��N�xG<z�f	 4�h��<a6@W�`��fഠ	N��OL{%rj��ue!����Y�1Ј�mwW1�	���8�~�� C5��g��l�{������إta�#s\ّ�?+_iI�!\M��	�����C��«��a�D�)�#��l S$$N�zO�7<ϣe�B�s�Ǖ���\�=A�`.[z"���%��{
�+���q�1)zt:Ȇ��j����S��9t6<��$p��Ѓ;��5����3�QF�9N�$s�y��e��x�.�<�tl?RwT5Λ�fzё5� �1�k1|��?Z}���ܪ'v���͈k@> <�$�F`FN�����p ׺j���3��
^E�?�}��ġ[�A�>�t��<	�����-3�=��7���[p�,�����h�Ħ����e�a �j�R)i��8�<{c���-S�*��s��J�$ �g�v���l_w�.KF����/��N�;����l�5�㈐�:�*+0��O-�8�~�����
��K�ŀ�����5�b�$�ʦg��,HO߶�?-s'1b��LB]��j��n�6�7�|	[�<P"\ў���~��BR_��U$ɫأ\�غF�!p�x��(
��jz�s_�%Y�A�7�u�?_����>��`���"��خ`�_�Fݍ�[[�t�zPK�)G��"��`�ft3�Z��|�o5oa�_\����d�����#5L),K�Ip#jaX�
B�_���i��
�	d����H��a�1��^��2���[Xpj>�_���?F6ܠ��xO��)\=r�Uo<u�S̔���	�i��.O��"�ɲ3E
S�	kqKV���⢋C/��H;l���Z�;�EO��P]XX	ތ�hf&}Ll{A���c���G�q�c$�}��t���r�]�<m=��e�K��If�j@������m���7�_�c�ޏ����z]a,�v+�:�9��Φ��I�av�������b2P��Fj�7/�h≫f�Nf�*��:X�<�m���r髧!-�A�C�j~?��<rﴶ����l+&3�>�z{ӽ�"�%ZFg� #�R�	Jx���_�T�ϑW��Ē[�;-E�בM��'>��bS�<N�qi M拯�\��+���D���"`��M�N1 ����3w(�[���,j�7�����C�����
g��3$ec����e�N�$\�@J@̖~�#�Fz�~����L����� �49V�������8��=�F5��K�:u��,~6��.}���R��jTS��\�R(5&l�G�C�����U���
����VT$�q}����4=u�UA���v�n���7��#Q�v��׸�T��fц�a�)��Z���%�۫՝@�"�X�gЂѻ#�0�ˉ��6��}�X|⥊�s��9N�ݯd��-��	(�����e����P�<�R©�z�h1r_�(Ak�l��RE��Pͺ��a���p^��Y$�W�!�]תA��ʴ_��L5�Zn6sAB�A·��*a2�͒�����7,Jf��~"є@��U�C��`�Z�g �Q�)?�%$r�zښ���n9{rj�r�T$I����!|u�-�pN��}G ��V��E�._�E��<���1# ��ذ�n�7v�E�!��u�v�Y5�_}�6ի3ѳW��*M��UF���5n���W��H�=�&��|/�d��tD��ـRE]�°���'(UUē�M��;�8��7��c�ߍ/H�_�+3���˲?L�`�PO����Z�RI5�XI,�ζ�Y�IP<��&�b%y~�����w�ǘ����4��۫4DY�M���i��K�ő��I�&Y�:L�>�n�)	Z���T8�����f,"B w�s�@�u��-t��	'���|.��F��!���F!;���R�$��CO�kQ�;������?!��&dH,���|��٦\j*�0�C��j��H>W�~�Ǣӏq�2EJΡ���s ��?��]�K��(���3�Y����ѐH�4vv:�f����Ъ��:���oc.8�����ٵ��k�p� f�V��ur��Ƒ5�=��";���J�(��s)D
�.�G�S�d���U��v�2.p�	�F�T�-f_aQ�[����f� a��a<y��榡O�U�aPG�Y~�cO[�.Ǖ�i�{Wb�@��E�0J�c�g�R��(�F����M�p T���:�w�L�����ܗ��:��7�n}�X^�'� o�gf���T��N�:�0�O�NNj屾.�!oF��pe}κ���j�W�j�S�s�I�=�o�R��2�S���]�BfU�k@#q]��פ��A�d�h3��1L-�2T��.@�}N\��vg8H����=���s�
��Nc���%K���Mۯ��Q���U�{���c��^'"\N�0ӳ�M����`�N����Ot�-��EN��~ߤ���߻�����+��~��OG-��E�+oSG��s�/���I��>�����#ƙ!2��cs�낇�.�ވctcW4b����Y6:A��FXAp3�t 3m+|����RI��.��Se��hwQ����A�#v��r)��9J:{�S�&)��|�3�[��_� [�j�{+:-���[����-��2�3�:�Gԩ�z�(�QT� ��5�|��ܣ�����/!5I�O%�Lxf��J4�]��ZSeo��7mبq�8	�����x�e�
��oX�jS,�
��_���)�W(6V�+��/�����о�>AH1梗J���?�V׋ �T�)�w���Ń-�}���p������CjֺI�`��.� �)�W2�d�㱳D��\�e���_d�x�sKET�5���q���؅����zY'm��'Uc�)o��ɗ��ׇN��"�:Y��f68y~�鯱������A��'꿺	1�O��&6�x���i7@��9�t;��'m����"R�w"�P��&�w��7^�Ϙ�t��� �F
^	.���nV�Wf89�+OYԚT��-��hfq�M���h�X��9�h�M���m���2�U&��W��!���������Gך�t�@x�͑���tS�e,��'��j���%ݒn���s�B*�*��'jaN�!X:�O'��$Eݽ#
��:=h�OŖ�c:����0��r�@��j`~`��C;�j� fc���`��ؑG��\��`) ��b���ww)"���n�w���!��>�
7C̚�Ճ��N��l�� �\0�w�#�׭����@���X�1��V$1�F�;����x-�(f�#omDc;2��L�BG����՞�����	(SY����m�k��ӏ�-���v'�5C�V���[ӌ�����5A0�����(j��Yƹ �k�Q��X�{�3�N=h"���M�t
���Rbx�IPޛ
��ޛ#b �����M4*�)�|9j��.��+��7��wO�wƙ�^�]x��)�C#�J���ջE�%�?p$h�z���롢�K�L�wqR�v� Hx5�����ll ��_��'��P�	*��o��Ԫv�����MOj�"�gcl�1/.F����bL�k�p��ݨ%|׽���sg� jj�8"�h�-��c�t���WQ���W0�xV�GUe�q�����v2�{��2��u�	��&Hŭ�vQ&d�:���n�v�#�#�������,�Ͼ, �0����v2\d`:�%ʚ���nw
��:�Mn�����8���[���%�D�������],�$�(՚]����6]
Μ5GF��Wr��Wv���S��vxd��(��o;9���Ӱ��Mb�=�nM_[,H�ym��?ɸ�����(J�⢟d�3"/�����>��6������b+�G�h�s�����QY�3*%}M*�n]�&���uX�/ ��_��7��q��Y/��ޕ���������S�m����t��nc�ф�X�.#�����aʷ�RΨ�Q���\�����6�ũ*q�EC0H�A�p�A�|�8���j��ˤ��Վd� ~��B��o���gm�-}���$ q/�yݧ;�9+P��C�ˎa�� {�*v�dD�{���~n��aU@�O���ů"���:Ƀ��L�_�iT_�W'}Є�K݃��5ߒ��hp�~�·ѿ�\�K�"tS��/4�ø�����+����hȨ�k5�*�P�c��QC�̏���?lE��n$Q:X�YA�[<?!/Jh�,g���o�}q��&�����c���h����i��6k����V��W	�k���G���DA����-��~��^y��1��F�Nz0&�����nՋؗ�"/�L@���ȋ_엘���>��R{!B��֬�*87�O����飂��-�،h��`ڥ���$�EH��I��(�r�lt�B���	�z��<#~8��������έG��vX�0[���U��l�1�G]�	t��iF��!rv��*�=wyg�
'];�m�&
{rc�R� &�"����ql���)��x{ԇ���(�B���4YǄ�9Ը!��JM�`㘇`��A^��d.��m���B��u�����)�JRk=��o�_���)����Jsz��j'�R�R���R��k\����|Ɂ���{�)pJg.j�J���ev��5�����J���+Н`�dfQ_ث�!Lo%�mY��Z��K�T��\]�H��a+R����k�vī
܏��d���쒪E��}����̍�"�x6���~��zm�JS����ːu� ����-g�3�rd�$7�c��5&<Ľ1�η}e��ay�	(�&��A~���2I��/��o��`A���<]�0����i�*�l�AL��D��/��������X�Q�[H�"���3�a鐩
��fxq���qO����Ji��4�4���S�<qh��I7i��m�}��7eR=P}q'���Ҕ�cxF��uT�� J�wU"���L'S����_ټ�{�"���>02W�K[��bSpm0�h��#�T+����;��Ro	u��8y��L�c��}8�V�N��y1�8�$BC����'Z�h;=�T6I��mB�v��):`q��@U=_�Ib��Pbjw�C�v(��Sa6���� {S��Ξ�_��vY��7 T�X�y1c�U�M>#3�2=���m,VAC�	�����9K��Z� �ŝ�[�1J�ԚUi�����|+��ͷ��<Fv]M��tR{����c*�8m;� �����x�⳱)����>�[�*�Yn~R7s�	\5����~vȺHi�V� 6I4Y��`�F��z&�x����z���%3�.эj�f�o������dіx���`��W��W���C�N�6U�
�{�aλM��W��5����5i�KEi>�^#�L�R9U��LwCQ��@(f�W�rQ3���������x�P��򓳝�}c�~�	Zfr�]S�t���W��ǯ�}\��+.k�Z3<8�LR=e�w��*���K�m��;���͢ۑ�X��+�Γ��L ��2z�R����V��X?��YGG�a`�mĬ57Y���MxS�޺�Y�Qy+������^.��[�[;�
)^*ß fq�#T�W��K��_!;�|Loo֘�o��,�}"�ͨػRn+� 6������A�X��5�R�-R�D�����U)�ظ#��{�(��	I��׏��N��vu���M�����%8�pm'^�'��b����LcJ�O�m�1��!�k3(A=�� m�2�U�[79 ��o24h )���Fa�4��.f7e΍K`�"�,��Y��1���߁�I�,q3짩3*�?��� ۻ�@�c	jV���i:S��B�̭o	�g�Ts'�H��V��3�d�Hd[׎sǑ��&o�B��I�Z0W��*�7���+�aU ���)�Ns��E�,�?������2��S��2�͛9T�Fz�.�_�G��>�
����/�@�7��.f)K�g����*&�ķE�6�� 7$����7Eܧ�� �*\�J�V�J����}���K�j(�p�!�j��?Sk����-�%�`'�]����ᓎ�E�!p�+-����S��Q$����������W�� #v�*Җ.�Qg~��2A[%ͽN�mC�h��C��s&���a���V�~�fc���9�!l#�O���9�-�i��)ƹ㿔���eoY���^�'Ir������U��T5��1 �K�֏�Z<oL�����y~3sf�5���ڟ�ߩд`Po��"�|�27��&sTC)�'�g�N^|)),����9��Jҷ_y�p`|�)�ױC����X�my�a�[z�������Z�Vབྷ!a��F��}`����}C.'b�l�������h��F ZX	 �m�ۃe���1�k����|�2�1���+#���9�/�
	�}���)yɓ�,i��}a�ǿ�V��[����Pk�Wu�Z��CZ�e-WAߟ���(��mw0�hP�U���?SnI��5�K�s�GC��ecC��f�(x��TVŌ��:��<�)�n��� %#�˻�f9�A2]��cxỆ�ާܝ-<@Y]z���Y"��ʠ$��}��\��f���~G�ƊNۏ�tw��#	S	����_J���n���}ۨ��c�ک�����ɪ�ɆGB�;��H�U��9����r�~U�"I"���|z�`H(۝�Ukf���4_Ӓ�·�&�a؝��G����A���O܆�8Ol'܅{� ���R�?�V�����΢��=��/96zgw�~��0<���$<��K([�����]�k��rT�.�}��;
�=ɋYc*�ݭgE���M!A��q�,�Ѷ���ʴ
7X�r��vզl4ÞI���_�������t��
�牯g�J��V��i�
->q�����G�Ĩ��ޕ���r/�c@�@f�9�����g�����˥	m�hA�6k@濼�=��s(PP�q�yh��Fo��<�;?�rJ,����l�!��E�w��}Z)P��`�$E��5��O�ݠo5��F�}Yu��z`����f���x���M��X=Xq��)Bf.`-?�g���<�U��(9.��$v�3��_�)ȴ��Q�ݍp��jiON�6���#���������.���
^�YDKn>�������H��&�B��'ܸ%e-��|�lގs�ɚ&L�$ˉ���[�I�F�"рr��,˚p
�P��r��?m�.�@��!NDkoi���N��%��h�Tp�>#�Ӕ��{��˂��f'������l+�cS�@պ�S�h�Ȋn"��|�k�;SN@ۘ
I7<f�:�*�u�3X:Od>���%Pg�A�h�U>Б���Q�T���g�=%
�i���R�E��+/�*��S/����g�~شL�4��%�A���#�x��'UB�]�:�t{4j�ľ�?�ΥD�BH�駅L�#�D���aK�6�:�9kFX��obwy�ݐ�hT�,�A���Xf��2B���L�K5�T\�3h]R�?ª� ��t��K)sF~��j��'=�(��W��**�c.{A`LD㗾�;(�h���;{�g��x��J��xz�*�T�ʣ�|��
�ģ��3c�4"�v��4BU-q>�>ȁ,Zc�٬�3��xs��dV�*U l�H�K�J ����u�Pe������I9��&�b����.?7,0���%��^k�a��P�? Ca��~��.��1�dn��oA���ߛ4�>Ӊ�p+W�&�$��~o!)�UR��Dg3xZ|�~�
Z�����d'�u3�	�W-R�\>� A��u�"ؐg;N���?��œ�/؀�i��|����\z\�hc�c.�I"'���4�j�d�W�nɇ����]\+O�9 s��jQ�J���V�RNn��'�)�AAK����'!#C�У	��������b}|�>�ƌ@H>#љkL���Ȧ�J�n ��=+�ŏ��&�_�&?I�v�\�Z��(��ЗT���{t�$������(K�P�\S)�x��ѭ����é��zHĨ�S�b��;owD��i1`e�����5�aJX�4��~x��5Tƥ.�����W8j퟉�@�B�\V$��w�L��~��xG<��-�5tS�`�&=�޸�����,u����Jפ�a���V���2f?>��Ϻ)0����'4��|p𰄄��|n'f��Qf���~|U7�#��)�����?�ϟ�7�g�g�䑲��ԧ|DmT����CUn��7�Q2�?� /���}�*]Mkt����ފ6� K!U���l��i�;z�_��d�������8����)"`�}F���2ݿt��e3��Z���yedͽB�m㰐L�G�D����v������E���M�����4�q����.\��i���T�j���|(,�|Պ� ��8is���c^�&��'NTtaX)Q�� ao�zE�`85ٞ�%v�$K���w�!�C�pO�)���T%B�Ŝ�����Sڟ� 3��s�U=565q�aj�W�i׺Ku�I��X��K���p%��W��2�ëB|������΂�d���l�5x����R�՘_Ym�Z�z~�p<���US-`�'Pj:x�Eer�|C��!�"(��n�kX�ۢ�l��U*<�.8�qb�:�R�C[V2���D�a+!�o��B ���xD�h�&lƪ�*,ƞP��` ���Ǎ�Y͙gwROm9L)��Y��Dh�ET(���g�������=����a�A5$�ڪ`;_�Ji\u�0m�6n)�y��B�$����Wv��S����3�Hq�r�v,�eF�z����ª7+��V��*w�˱�'>��[0yVdu{��*ͧ�jX�H�'�����q`��c%����H0�jY.��Z1�>t`P�	9�1}%fb[Q�^��tϻd���eG�[
�A1���B$�W�=J����>��e	�9˴�6#zL~v���۴P��k��Jh�!�����;!A!e�S'�P��4�{I��N�q��'D\�2)�6���e?@/}�
	����Ьz1��	V��SQ�:V/6g�r��trf�O�`T�%x3}�$\�J��������Vv3=]�&1]���c���|&O��_�C�p$��{D����^�C�*L�5�`�m�I}�$b�Q�j,35�B&u�M�+�`�2��u� �f)w��/@�:�����VK��v���׸�J��4_��m�6��h���p�FƵЃI5�F�4��<���7f9� NQ�؏d�X�s��GF����5��ch�~ʲtO��\Vc�g�lTf�%���:�	�ƛ�h�>A�ɴ[����s ����V}���:���ë��M�?�_b�@9ӛ(4���0}kF
c���ļ�k=�-�o��K��Y����?h����c�Ϲ��U�$TS�^���?A͏�Zҝ����q3�̷pA������G�!�A0� ��U2�$�%-�+�����ʶ��*׊E���^��?���լ~���Q��!�����M�:���7�������u�NK8�S���~\�Yt �9��H(z�,�q9S?AGa� ���A��Xb��8�_�j4�W}v�E�f�p=E�F\G���}g��ٍ	��\fk�x���h�w���2~Yu��E�ֻ�����&B�P5/�4.F����J{�XD�m_a^�va�~km�k���	(���(��>f[7'�s�k9��k+X��R"����E�����s��I���%��*��j�3����A�������	��W�a�;? ���y�Z�m�l��I�/��T�����{"3<3.il�y��T��sp�`��qaF��v� ~��%��t�Q�SC�����rj0��`��L߀$Ah�=T��n��~��_DJc{���Aa��r��f���4t��66jx���;���.�F�m�b�G��lZC`��Ŋ��#�s��n^�ﳑc���+`��{��X�t�0@0ϳ`@� ��D���"��u�ž�T�?�ߔ-�&��4A+S������ǿo����ۏ�����n \~��	��`�H��t��a�y�} ����};r��ȋ�Y-k;�L����l�:5~�C?�8��r7\��m^5y�@��tj#xލ��� ���~�E<4�Xt������ ���@Ɇv��U�.֟з�1bd�n� ���YHT5H���j�.��h]�D�"Iݢb�8w(���&b�FJ��y.��]�49��vJ12<����k���gԖ:�;�9��F�R�a�?�ڠ1\�?ꇁ�����iq�Ѷm���@-���)>%QEe����̊׿yuA-��+j����loV�9B��U'�R�6�'�E����&������_n*5#�ذ�.��)�H����3.���Ky�3ڒ]^�!��]OJ������ʹ�m	��w�
��4oʣ�x<�����)�Ia�L�e"��De��SL%�����tB�	x_��8~���ꠦ4Ց� H�DƽK����4V���Q�Pܩ�d���t{@��Ri<Wy
s�7���	]�[Pp�֔º�c��v
��M�<�"�ge"�:S�*��=�D,�z�	��^���0�alIYb��V_����+t�3��߁h��)�b�������(:��x:�@���S&����~t�r�p�/ِ�H���(r{�uăZ�J�Q��d�y��[��zC���O��p��:����c�7�BA�.��YB�m, ��AF)�x���+a+q	;�1[�.'|{L��Ƶ�IXɡ�vo<����������I��?6�1�OG�`n@ \-R�$�w��ah��[�֭��9mZ��
Z��,4	u�1�0  �@^v�[����LeZ�{ML<s�y��/ؤ���3\�Kv}y�cZ|kY�t���н?��'.X�l	�YE��^��v�rdʪ/�F��'�6������;�C`��	b�O�9݃tO9��+i=�t"M�t��ǜ�<S��n�\K~ڈBpF�t��g���;�͝�KzV�;�}EP���A���,��N����$����gb��w�%�U�1H�Ŵ���Ԑ,̔���b7�[T0 p��D�/���?�r8�tq�z@����uN�OpBA��6�ߛ%�(E,q��\��$Ga=��lc�Q�	"4%1@ ���%v|���������I��n̈́h�8:��0�;��xv��	�ͫr�]9���\Vbi���ۯ޶�(@�2�m�4q8��[�P��
 ���9��ص�-r�����Mx��m��[��V���7�JB�K�݀�@���!��1�������]M�z���p���ѫ��ޛerR�[PT!��W��¸Q"g(�I��%�A��N2���e�F`��7;�ZK˨¬[B���X����p�|�#{������&hQ�j�P��-<}N��#�E!�\I�ET�t؅ 6B�g���yX����/"Ԭd�{}�S͠\uUcǣR�\�<!��̼�:$�E��BskZ׏?���C�yo^����{4�>��\ʐC+��A����Ԑ�up�1	��;��O<�}ۂ��z�?k	0t>�7ב�_�q���IF���s�T�8>g���ڞH: ��HR���`�y �{#jw���ˎ�ҹ������['b�y�����W�n�mv�B�v�5de(��.�hs���J�C�}�Ro�%��0��r��"ʜF�4U�P���p*O��p�B� ���0%H3��J�b��A�GG,��+q�Urd�*w�&��w��t9HM� ,c*��{��N��&(���"��FYn�EټÉ���#��H��� �⒈��2����e/�?�SsQP`��ʥv!��g�<��� +lf�>{|�a��n��9��S�	�L*{���[�od��c�K���3��w�͝�F�%��!V��![�Ȋ�����E��(;eZ2���6/�tM��0�|�
i���y_mV"��)�ֺ2P�A�8ޢ�[-'fv\���.��/�1�k�4c#<L�P�@��q�O�>����p(2׮�S_>�rC�����F��!�=:^C&�*��n"-Ͳy�WiQ��u�o�]+yF�����ȵ��zu�}����I:P7u6.޵z��ᛈ�urS���S�d�[U\�HSMi�B����t���P��X/��)����ɯQ9+q���[�O�(��yfҞ����'�Y|;nJ�:01���r~*pn),V�3�A�s�y둘m�9]B��Qs�@].�<����#�����Cx�͹�w4S&
m����������|�b#O����O���Y�Pf��7��+�"(ʺ�LƏ!0�/}i�>�1j[nT?��I�"$�cp�˻x�:�M�.���2���5�6���Qk�4;��KV�����T�E CJ�3
�yB D{��Rp�&=�7�8��'_�_���F	�l�a�oY[6��S�/��z��w��l�F�Օ�R���<����!k�<�dh)��$>��j79VDh�m���N2v
}��Ȧ5�ǜ	�G�7O�0H8ʯ乭i~��4/΋�պ�t�F��t����ӝ���3��;��x�6����]�ޮ��i�*�w3����4QT���Đ��T����J����WE�a*�z�2�	��l����.U�M�V� zO�ŨY֦S��.{G^W`������ʓ�I-�����~� ��,2G���2'C���J��z�M��zL�B�4��=�����~G���G�]A�޷�Oo,�`]����|�hp�R��%�� e��Gs�]���"b��pfy��ug�)���N�+� �Eu�f�_�8}=l���C�oD�{�dc�;\ڦ�-tx{�Q�����_��v���Gg�U%VQ+d6�m�ܧJ �d�t�_�-�Z���9"�D�W/jN�=M�]c=���:� ��{B�E(z��h"��V�ɻ�p@��i�W�£�.��\O�l��%B��sI���!Q)��h+Էt� yC��-�7��V�F�*��Y�����2��c����r?�	���x.]<�~��^�	!�8>M2<Hソ��鄭�[�;n����F��@��O��ԨaN���Q����Ҷ`��1Ew(��g��!D�ٍ�H�s!ޗ/��V�{�۵�T���5��qzv�U�*�D�SO=:��H
e�������kZ��SPs�H1S��M~�o9��)Bvm��
�s?��'���_�.։ �C�[abtJP��r`�ي��ў��ޏZC�v�ǼS�K7��J��)�|L�;4����Q0�fF����l�1����:#��9��wlQLy�:�yȗ�Ȍ�����x�%R?���TȽ&T��ee�6�J��U�Ç��M�� '�����p
��X�̾��]r�-�7����5�B���Ѡypn���1О��a硋��K�(X[�]��l�b�H[��C+�Q������i����x}���(�CP��~�z�����CЦEw.HO�]�ȫ�=8�I+Q{�a�%��M�<rΝ��W�yOM�+�w�X3�i��4L-f��@�@YF{J[:�Ix�J� Wߧ��_\χ��9^8��PD���k�M��D���bS �F�$��.u�׹ŷ�&.�`i��K����C+\�=�ƺe���r�A!c������}ME#�{KVwI���i,T8Ѿ3�^�1�§W��a�`Τ�vz�nY)�sOY曘�[,�̕����~Z�ײ��'%���y�L~O���-ָ̂c�@�dݠ&#ۋ�᪡�sa���!���݅t�����j9toAS.;�a�(d��1���A���ڨm�Q��@Nͦ5i�j*+I�I|�;"���C���O����2|�G:,�������#YsP	�ۤ Dc_.w��?	Qf���V�bR�����F_�-�?���,��=p�n 8h,�iq-�?I�K�:ڧNV>�C��{�4*%�c�E��p�\�0���,!��j��T�s��j�R�q�/�$a�N	��:Ǚ�ɠ��d�U+	:�Ԡ�41��ح.A��ps��(�Gl��i�k��~�`��[��
�����f�E��xY�nqz>[a�5�1(��xw"��ZL��#hb�M��1@��'v�64�w4���#���^;L�X��!�����s]H.h=o��*%��6e��Qe���jP �H��>��&��=�펥�0(�3��VT����l�U*� ��Ky�+�б7���1��i��H��S�l��i���S
�w^r#[z�ʑܢe,T@~CAӦ)��	�H�v��E�)b�I
��T�� ǈ+d��E9��X�ꛈzڀ�'����R� �a2U�m��t�5ݷ?|���p-�I7� ��D��X�g�ۨ]�\�t8罾�茞 "V�*�e�]��P��MTf6j�JRѳ�$&^W|i�z�@U�4���@Hp�9��M5n��v���肠#��"����y+!�gv{��cv،̎�3淖���H~Ka�oW�˚^04��=�0ű�<#�c�a����B�;�2�=���zz��^88��7lԗM�K���)�,��IFK�/+�fS� �G��޽^����t�:�6 �$�y.��mUJ
��H���%��G���o�p�k��|��$�e�W�ڨ���8��,���Ա_���@E��W!�
fV��SŜ�^z�9�����Ҧ[N(�s�W���;H�1��"���jth|��jn2`$�z�h� [GW��і�f��Ѓ��L2	��h���,U��@؊��}*���5���s��P#U��\TϩT'��5:9�ƈ�.Z�=�-���_
P)te@����*h�K�Lmdi �����A���3}PK���LU����4�͡������:��4��""�-Z��\T5}`�-ro�r�(AW��ζN��-�2�#�T��j��0Iyf�������H�j��ME�Fʡ�f#�Ph8���y ��u2A��I"T)�|�m�NC�4�vp�T�+Ћ�;@jB��aP<nX:�������Š���G�����9�t��KĘ`7��؇M�d;��	��SGWک��@���zɣ��.ġ �ԨT�͟��'Ǜ7�a46��b��p��� �=���%�a���o�6���M����\s��$|[�܂<��׼�QId�.�[[�L���w�ʨ�5��2'�o�`$�c�C2�p�3i'�[�S9�Z�y�b�����ۭ6�2��~��	�0�(�@�T���zS���;D���hV����L���\���o��_�$�>��P�$��h��Ǭ����*��z^O��x�o���;-�V�rXd��j/�<�0>ydL[pzb�g��o~:�C�0�<�����҂���vʳ��n&����C�$1X�	�-�?6`�x}75�>����?�>��v�؆ߚ3N)e��z�m���z�+'��$l���E����o�R��"qeҤa�`��P�%Yh8��a&Y�/������?�D��z�<����� ��d#r5���]&��v����ԉ�o��쓸���E!�Y��%���l��Z4Ąs8��Z��5��g<��zN3�D�M����ya)�:���ih#(Xek��b��K�Y��|+������ I�_DgG"*��͚*����`g�ǂ�g;o@ŧϕ���'vQj,�TqSi+2#�_	���H��P�Ȍt�.��T��{V�8@��G|��|��Rԫ�~ ���FC�Sl\�u!�9��k�;���-)��z�q�� FC������va���TIK_��� ���j�$���t-ϊ���\��
���Kr�
���Q�����(<��vm��BM�d�aX���I�JUm�H�ϗ-`1�s�� Zb��8OGHW�Ǭ���Ȅ_W��0t�,�j�>{�c=�����fk�g��G�_�[}�mK���T.�Sp�||���IE��K�E�OX�C��ϲ#x/c�~W��N�)��V�WS�fT���3h�)y�Ϣ���}ҟQG���O|L���a=T�z��8<6m�����>L��V_0�) ���E�d�V�4�\-D����&,��q��H�3'�Y�ȡ���	
�Y�H���Q�U6Pr�d 8{k*d:�6���i���w2��+.�X'a�t�g���:�Y�F�6g	�:�.�gP�'~�x�͛�?c�-}�x�m�'j�s�����W^��K��
����c�{,O27��9[�[zk-t%'�� �{o�Zۃ��2/����&�, =)���$�[2�:��)��j�ue��!�>o�f@�Ӑ�@����Z.�;��l|���_���BM"�#����-c�1����̸��y���W�I	Ӣw	�aJr����Y��ˆD6�o�Y�q�=�ږ	���d4�Z�A���Ⱦ����A�4�|^&�]�#J'T� m�U ̤��L�~.?B�:P���:��C�!rc�w�]|�������'��ܥJ�|��/���d�$AJ��đ�l �	+�����E#~K'n�<�G~�Jeμ�{����}��~-����a-"�.���Vp�a����<->!։����Ut<����BtI�`pH���N0�E�mu��`0���>�U�1�&"���.��e��Hk;�L�Ж�t��J:@8�;�lh�뫬�Hڮyc���B�˕@zU)�y�l��5��կ4�͈T��>�,y��&�#'�Z����X�jvm䈩tX�*L���E�t&v�7c�(�%����"Ģ����M�G1-Ϡ�=c�ܸ�{�r�T����J�?����?$�x��6���}nC��H�����\pg��e�)j�����&��vEk���]�*,R���K��d*P�����F��`}��Xm$>��d(����:P@oam�N4�M�ڛ��#�����꺂-�K�U�cE�O�bO(�{@�j����)E���&uL�S�Ql�g������}8��t	�O=���fl��[������k(��5Cѕ���x�Ϡ�9��\!��Raш|0��6�[B����IA�0B�3�E�$��U��i�[ӹ<}L�����<Ʋ�)c�5�_���1���n��gZ���g~�"hb�G��9NG_�I&����k=w���+�:X1鿌�<��W���u�zYh��y�p��(>�U�^�b_�ho� Sk�mm~a�8H�e𣔉�j�K����yw��r��Б�X��p�9~�-���UiZ��g�[�O '�ĩFV�4�� �z[��{C2���܃�\�ǎɠ��m���3�+�ZJ�&̃�<biu�/� ݁ �]�tSUb%�ƶ�+E�Q��<��0܏�F�~X32l}T�$}���Ɠ��� B�adTx(NrIQaAĄ&z-��B� �����2IP����EЂ�r��+·���e��K�9���YT����5]��An0��{�^�=Z V��N��g�B�%|��7/���m(���%f��q7%��"!��8~�?�@�4^o-�X�k��� ���E�aI��»��,�B��(Y��t螟P\�˰o��I�FG�t0)�s�Ge;0�w���jgxb�j���i����,s��7�U�$ǅtٳ��<�W-��GP�YÞv�H�:|4�}���+�ŒE�h�\	c5\0ܮ��|5q���g��
o�Z��ΎeWV���Ӳsri^8ɬ�۔�d�a����jW�  춹fVmDQ�m��N�!HQ�T�P�>����\:�K�$:}�74�[�V�"��-�4�?4��1�p��ފC�1���b	|&�̚9��}4OXaJF9���ѮSg�p�J|���7�fI� �L}�d�Xn�E��H�*=�l�^5��e�iVL���X�V��N�:�e8.u7~Xx-���,2�T��D����y�ӕ����h1����G�?�KqBE�x�)��k����_�97����+�۵�W��5�|��x~�-S��ԅwߢÍ��ڨ�A��c�%��m(t`&}_����J���af 9�#�:�;L��b�ȯ=.Qi�t/<"";PXD1����Ƥ&[5�r����@,���q��%r�?�ߚ����U��3������1��@(����8oZȘ�G`�bp��t��6�5`�N�<��#.��O��#��ω�5�=�u��&TGд��W&�w���
9(8��,���LDo_}��`\�U@a4^������tKX��P����1\����#��� �ݞIJB�1�m���ҔI\����ع�Yر��tE�FpD9D���6�M�A�t��@iM��?Xܟk��u�����ꏻh�OaV������Z�L�� �}V�L'G��y��(A�j�R,�ppc�j�d�㿻��.�Ag9]����Z��M8�@_�T���=%��S����Z<�Kc�ʲr ��Z�Ҽ�f�����J�V5�u\	iAPln��Z,K!ifr+ �'��J��F��S0�	/}� �1�R����
V�!���Q�@ܺ$~���Q�mBRP���VO�NW���JG^�J�>�HG�H�	�H\�l*È��RW�G�g�Ye�Է��K�Y5iG)�B������1��M_�H�BRA��S|&��9��ڏs�X����v=�O5�FXp2;�^���M��,�*�#�RMuV�-�؊yyLH����cF��ᔚB��C:fǕ�гo/Q�[Y��h��f7�1�5��K�v���.(�N�J2{)��!{��0�M���R8�yda�N�}R��Ê��%�r>?A�A���l7��s֊��F�1/m/H�|'�jC>�����ݿ5������^c���BW9;J��; ݱ��V}�X�R)h�f/s�;�����8$�����Z�����@,5�!���>�"��(Q�e��e�kUZQ�N=�Scg=�ϴt�Z�=Dwn���q>8�臚�1N7���=�N'��D\~0�X�/��Q{r�o��|T
ZJK`�����+��:ܱ�Q%`�p4|Nbb%sG�f���:�;�l@_����Lcث֞�B\@��c�E��~>u:�ZN�.��Ƥ�� �A�r.��-ypVE��Ee��C��(�zt����&�}���Tp�Dn���׿ꃼ��&���2��d̀�d-M�Ɏ�0��S\�^�P4,Ċ]�{�m���?Ԍ��h���ibɧmP�ޡŧ��{K
r���^H��F�RKU�'W�7���_�2˫Ñ JNLi���"鷪h�z���AW�;�C���P�n�d��,_� 
�Iw+j���� ��E&�0�  % �$u1M��0�%��E��dy�-�7q�2m�Ę"�W��묓����<��U�w�3.\�@X�2CGN ���[zY�?�u�T���MR�M���M�G`�t�u%_p�E���l
��)���*&�+���YK2l�'J��2����.@%��h�y�0�qx�٬��VX��t0<�hp����I4*��0�/�X�h����K�E���1�{%�P-Ůgґ4D(9���%zZ����j�$wm�b�z��� Q����O�M���U�q��mqC�D����Z�R>�a/��1K�\5�2_����q�V	��c� �/H���f�h-�I��1�܋#'nm=&A��2S�JL0 B�A�_Y4��n��ۺD��@B�8<j��!�Kj{z�ǠJ�+�귐S���i�HN�T@�n��Ƶh�++�/��HN�Dx�~� �3I��\𬞏v"��*�~ӢG�j�߄�f*Ԃ�M)�n��^��ۿn�4�)Y+��|$�EMz^,�w�o���HAɹbU �̋%�M��!N�d�܀n������5	�)�m�Vi#�w[�b�RaHiu/�l�[��'>Л_��g����!!��N�(S�Y\˚B�0�t09��D�kv~��3^ȧ��)ux�WfSu�p$YW�U���'�t���~ :�7d����xj��W7d�Ƞ�v����izi]yn4���9E[�Tt���z�*'�Q���s� �ly�RY��Ś�m�R����0�]C?�C^,dp�.t��.��%�J`}�Y��Gw	i���f����v�%P��x7�<�Y�%��l5�Wcf#�2�ܤF��#3N�Msi6��c�^ɚ��J8��� >=��= �h�5C�yMM	\�2,��+�/j����
��5�;�	o�L0�,0԰��"[�-�rJb���R�큟c5{n�<#˷�ǚ�j� �h3��Y���Y�y#7����y�sԀ!gC�ƥN��[3�kBl���L��V��ӵ��l@�̴Y
r|@�B�^JI��-P�$����%9~��������;���+f��V[�[��AJ�bǉ��9&)�Y�-�����O[���e���j�[*g�zz���Q,r��.3�� $�N�ڢ�˅����@P�H����� ���3=Z�Y��敤b�v��u2���`��'i�>��w}�F�<��\����:�k'ʜ|����KB:Mum	H_��]�H®}���@g�L�Z�i�8v�	v���{_ ����+m�[+�W4`� �:�EB�"���~bc.��/��ǧy��e�K�|@��p��k�p���ld���E�6X��,��~�J��<��t��` R?�< �m���ցb�QE�"���*�5i��jz5eߗ�{�TJP��*�(�8*!���}jn���K��
��m������D3���Y����pPLa3����ԕ�0a�?T��u�M�>{�^�@mx���|"�"�h����Lc�B���Ayd�=r���C��]�PB8">ď�JH�;��Ձ��i���l�NduK�RM؏36V��n��4u�5W{�\��z��2���o�T�@1T� #T���Q#)�k�)+�`1f�o�g���yy��י\2�B��¤p*8� ���=:j"��3��6
��a��i����e�A�����k��kL�$؉�y�#��`��S��}Ӈ?�Mw���Y�����dBy�!L�N��F��i�h�E�xqfL�N�R�3��kc�
��r\��>� �}�@�KNCrMoB�ޫ����!��7�5��N�k�V�[����òj�15:4��dnIfq�Pl�&D@dS���YH�R�3�T{:2��I�e�H
� Ą���9�g��ޮ�K�����Н�����'g}�QS㟤We��r �/��(�i��ST[-�S��P��q�5�)�n�ȵ`r �4ͽx �;FS՟ O��c��TK��I
������g�Л!l_�d�5�_�[�P��eb3�,@��
�ˑc`:-7T�@��S�p�l\&���cd��a���R����!�赐��,x���w��ӰEE��}�DU��e�3�w����G3�8��� ���c�(T����P�F=��ǚ�/
@P��G��-[��p�ay�W)れ��R	-M��q��F�Y�_�5�"�k�����o�C͆UwI�2�BXoTv
��8�>hwCX�@�+A5��@�`��y���K�9�oI�����.�n`
�*�����E19�_7�gӜ&����H�T�,���-�ͩΈ��ц���h�8�zDI?��~��p��)�;B=�����^�&��h�M��a!H��|z7�d���\�YJk��6�ġ3���-��ͻ>�l�{�Z �ǎ�Y�	lX{PAjU�h��<����?��.%@�m0�`�Ԅ�����ߞ|Bp��{�Mڶ�����܎T��!���^���>/m]���3		R�>J��(���_��\
�5�j�-7@�R�X��Ue���A�(g�2ԙ׎��v�q?�T�F���,��/�Oa �hr�p��� �B�v�l�4������ו�γ�|��%�s�w�94ڰ���8�V~��̳�Ci0���D����Ɏs�o�i���lH���e!�SPW��'Cw%p|z|�W��,{�������rU�����qr8~��W��f��;��|���C��19�/��R���A�� R+v����s���bv+l� g��xz���|j0r����ya��(���z�⥇.��ڑ��rua�W�L�1w���`�u�7�!3Y��/��KN�������8eA�����W���-�ϟ)�G,|��<bͯқ�g�C�-V�0*&�#���Nr�M��
q� �߭m`� ��j(������,-��͔��	��|ģBI�o���	��"��{d��pyD��g����p�;�#�N�g��s��0_nz��b���S|��[��|����G�pWQި����xk�	Y}�%�7JMg�f�c"流w�w���e�3�E���ײN��sR*�І�+�x�%�"Zz�b��$,	��x@��^��d��! �����޶�2��ֽ0�r|�O�L $��`�29׾]<|�N���D���yk;.߫22 WgC-��S�U���@�1��)p�ʻd�K]ܠ(k��6ٕ��=����/�������Ԣw,AmK��w�4w[���]v���+���Bg[E�]��W��x���(���Z���1cf�[�C�OO+�T#�⼤s#JY=��'eD�_�/(w�
X��8j�.EX{��ֺnWPaK�n9����|s�i�.:Uj� ��� ���"�;)��"�͕�)u�i�Ŵ��K#��T�Gmw.��|]wv�ڗѩ��˔��Y*n 7}K]�J��@�j�#g歿�lc��bsj5-�B���9����/��+��p+�Y�8wyE� ��v���{�^j�l�q���
��=������? thȘ5��A4�-�~��"9UZQ���B�ZL��Ԡf 4Oϔ=��\g#y��V��)�]5�C��3���6�jh��IU���$w����Q���2t��K4�Υ~�\Yߨ�����'����[�'�8p���Em��"�6������X��?���C(Թp�F�y����֖ٯJ8�U5���a�mH�u{����h��U�Z�Qn����vĦ��*��H�eC�˿v���/�� 3@���6F^\́Cۢ��%�*{��8���wLt�sRez1F���o/	�#а9b�9�@��sP>���`	�8�:;�8�T�<��Ӌ��#�@J}�T�t�%m�$���g4���j�����eJ$��zH���9��Hlo]�RMSA�G N�]x�Y)1n��G��d�.Z�|P�B����VFČ�#��a�8�_�-�SC�:Q��g��#,����ۀ���ئ�U�K@P}U&��?ύQCz�Z�������(-B[�.}b��=>;n���|N1�M����dK�G�-F>�e��G� ��:���^�^x�5�ڤ��5XI�H��=1�����s1n��8Ya��LM�+�P'���yɣ�m����������;��U��I�g����]�N7�>d�J՚sp�G���P
�@�F2t�����m�s��V�������C¹;�+�s�����]���5t��K�BL��e��1;��v�`���7���ȏ�SL�G$¡E�_j��\k�t���[���b�i^R�E�".Y���ϴ�k���7��$���=�Coߑ��s0ٔ�Z:VS4 ���KF�1$���B�v��q�0w�̰$I Ȩ���Ǻ�M,�QZ �I�Y`��ٗ*q&���j>��y}��G��������ws�Z!��{�i��K�1�U��/:L��b��Q�c?	�=�J/����3�?�w�[�SiٴʸÍ�JVh�F� �F2qvx�ۿ���Қ]ܕ��	/B�
�9��ҥ�ySH����q1�o��t�{���WM�\�x�_� *i�Z�~1_�&���X�B|�A&~-cS�M�2R�e���N-��`�>֚�U�0s%<�ը��ie\��9A7��V��}1�[KɈK�
�`�xY`��2'8���!�M�!*�3;P�2�ހ@M�T	���v�{"��b�q*�����[fAC��
���":��'ꪜ�>���IX��K�qrW" <v��c�sރ?��*�����'�^x���@J�B�yxe�)@�u����
�sE>5k���ߦ\�}l <s9���[���x�k� e��5/6�C��<[��\����ٚ�^��Bc���D�ʩW����
�AK�SU~�"���eL+e6!T�F�R=x�������A�KĔ�kIq�dL�\�hs�H���m�=�u<�F��)/�D�4��@����j�W���_��T��9�&k�M�75w�,�X�<	��9�ղ�;RU�|(f�ց5ha�l�^\��ڜ�vm".2N���2�|�u��&� ���u�	��7�亜�7ltݺ
��)������I(^�J�u#�� b�?9���yׅ/Y�?�Rp_5���W�4'0U�#�H�t�vW�f�$���I�<�ϝ��w�$I}
�^Q`%gD�A�-(�*���? &4�t)B5W���,����`nNG�y^@Pl#��d���=���	n n�o_S�do��.U�ԃ[B�<���ڎiG��wYEH�᫕�	�^����36^��b!���Y����^k��'��b�g�t��}���ْ�1�M�ޡ�)=e�i�?�E����2QV}S}쑄�tt)e�QU�F��sbK���Q�w�wU�<�pm�VX�(w���,9H�1"����^����X -�Z���u�|s�%�����QѴĐQ^�o�r�"	���a��;��z���H��E�p\b�4Խa�k(B�8_{e���n�.X��%.�ml�&-�~����A�7j�
�[I�4�K!����G<R~H����0���6C�L����`X�m�E������B���"������a1z ܽ>�{�l�e�����-���7q�A`I�fq�$	��j{�; ؏+�1`7�W_vS-@�	����F��/�QF? �v�i�U�y����$�;�H���B�l�|.+��i��\���h
�H H%�l$&A!�{��J��zv��:��r���b1T�6��թ(�%��籤��H�O�\_����l�T�3���dWF$"�0ɓg����%O�76;3�3��Tɪ�Co������S��I0ͽ����0�w$b��{g&j���NA\7��c��7�
���c��J�~0Ì��C���?n���j�r.^�?����=bb=�r��~WV�C^�����wx��
2xQ�O��vpO�:�xՓ�)Ξr��̎����!S"/�F��Ab>Q�*$�n�ZVKJ$����Ƚ[��My�#m|`AC������^2����V�?!��?��e�t
uCŲ��H��(�DWPٔ�����8�n�a\��7=P��B�ƿ2�K�_z�7	�v�6�iH�p�@nb��#��t�J�׮~��
�F�������%3�:ĳ=�R�g���C�����!�{��m�u���'KM�o�p5eRN��\�uz��Ԅ_ƿ� �i־|�1Y~���NxB/���}(���x#z�n�0ܤ��(P�|��;�D�ǳ�Q`�}��>�'��5'������U��'4�z� *��6��JoK�W�M�D|�x͙�#�"'�S.�0d�/���K��M��;�V0C#�����oB���{�q|9�Vt���o�y��G��*�5  wT�v�;f���{qf�E}3 Q y���f������e��FɅ\���N�Π�����gI �weAӭ��.ŏ��v;�/ş�ܒQ@Zz���z�����>X�9%��죓s� -X�y�V�Gߒ�=�>939�G������^d�h�K���[��LqW�D��O��L�fI��3��ocA� :0A�	���}��J��+�n2�������]�FY־)���$�;�@Ě;�}���	�RҲj���)�f�@J�n�r�(<����Rj�vv�~#Ǹ�4�1�4��ż/�V?�u%���nB�v����M{�W"f�T��ab��٥Du_j���k��u���1���0ER�vSʿ�ҥ[!�< T��U�w��Q�a!�F?{ �dW�	(�[��X�1����Z �`�Z��TF<�F��&1�2�NI�n}���E��t������Uܮ���Tg=8���J�ב�+[��ݫ���2A�I�9�*��wa{�U,�OX�|v�	����Om�l��AN/x|�@�#P_�[���%w0��ҦT�l���-quu���n�) �$}�Hp^>�bv�jڅ)�u�� L58f>v�ճW*/s[�v�=͍��NKv�l��/����Ak���
e9-�V�_����*Ā��\P�N�k3$�5�Ι#��$��(�'ٱ �=���t���\C�ߴT�o��N����-�׭gF,�(���D��?8�&��{]��cS��<���zxlƀ��j2�o�a���.��U|a�����������v1,_ȭ���x���D����9�ih`�#$�u�ĶI��V�<��b��5VLW �����=��	�� `�#ᷣVHj�5&�.�%h=�U)����P����I��^v����s�'^����f��#m�e�1�O�`�ꯒ��A@$}�c�3/"�U����J��N
��
����z��va;�1���:xYE��om����Z8Z�tA��x.� �F��g�����F��R����eT9@_PD�� F�p��H�tsZ+t\�� �0x�~� NwO-M��q�0h\g���0�O,�09p��:%����(HA�o�q��^��µ��YD9&d��M.�3�*"� �V-��j�3!*��{���V �.N�ɣ�o��Fw!���5�o��r�����:ʋi ���f��5�Q)��	�l��ů"K�:��B�z����Hg���3�AԶv�Q�hg�Zd
n�B�l�R��)r�U]찭�M��<;R�\s�0���I����������RK�}�X&��0������ �g���%�=�@Wu��%=o,��= �����^���Q'%O,��z�|v6��f�縊��˂̘Uq9�y�(��ݒ��fQ�Nj��� V��B+T�j�8�v���6�
���@�|w�v��A���gk崫�9���/5[{)���J�)�{�f�:��]ى�:�� �B2� ��cWp	LMw�q잳�@�:�ON�@:p��Ճ���^�:D4#[��R�x��1���y��?x���_�N� �j��:/J��Ƹ�qX�n�����G���r���P�F��`�X�FX[͵��ؚ�:�/Nr.�	H��ј;{u����ǲOo��WL�n�?�8+��V)��!��k3/	�d���<<1��3�����QY�S8
�x� Ug��EVׁ��S��
>j�ί���J��@���'M.�><	w�/�f�+���癅���(68`�'_Y]L�����`GY�!]���)~1$���U~}�Z�u����%��S�F�'� �����y��_N��e� u��a/� 녾�<"�+����Sԁ�����y~�`I�	���1�۽�?􋢇���M��4ٺv����x��������C���:s����u
�`�%�IEH�!f�V�C�(����(kS�'d�a�v���ݾ_RSQo�g޳+�$~ld�-���R�������$�5��h^�H�U� �4�Z/4
�)�}9�C�����~�3� p@֎b���}����`]x�;�X�`Q��Ǻ�9Q���9�%�JXP o+�MX�o��bfq�t<w��#y�
�"��ƋЙV&h��VL���g����H)/��I�
dp|�{I��R��#(ն�-����'=~�UeT2oe{̽R�!�� �c��8$��{�u^b��Ʉ�3�R��g	���p9ݤ��0�*��_�@P�;�n)�J�ʦ���������-��_ͱ��w�o���}�:r.$ S���h�]9r�R-t�B���K+�'H�S8�s�����O]m��_e`��]�P@<<9Q�
_OЭO��.��4��}����̪%7u3i�����9-��{�y1D��7�J饹j~���2ȡ�/���pg�tP#�-V��9#����B"�\��h����t*|������9�(����\_��,��^x� ����j3��z0ͭ��$�>2��9?�e�I����mf(B"
�!��(&Ƈ�ˇj�*���DY��*g��g�`�//�	�9`��֣�7��ң�N4]_vm�!@�2M����#�Y/�`����˛�!+�̲�3|���3F��6{0B��	��V����~g�g�`P/d�e��xZj��(TN�t�A&S��8���ﬡ��s
��ݶ)�l$W�α��L�ƸlQ'�4���	�y�m�Ŀs�߉��l�RK�o���vڛ�'<Q�䐉�J�I��N�
����r�>�����\�<ްT	�uo��씖-��p?c'��A��S�6� �f:5�q�Z)�_�l�0׳1oo�*|���2|�g�dU����q�� ��`+`��$��.(@�1���X~Ҹ�z��$��:!Ώ�V��''�IObM8_c�̈�̭����˨�E�oSp|�n��_y�H�8^)�g�!��=�0�H�0��N�kL� Iw 0��"�K�� ���l&�׾h_���[�#ܤ�i��_�!�K�qW��Gb�Ԡ�(e|(���Aq*Q���#h&��s�F|�x���a�|L:����ʂ��
8N���#Y��BRi�?B$���T?�,��f����L��y��`�sd
�- t�����!�h�8t�p(�a��|��3@�ܒW��P�Y.8�����]t���!�:��w&� �����J���:�E�Vc�����|n�D�Ġ7ǲe�V4�$��7�cC�3:\5,;�j��Mi~�ѩ����<I�EA�/ &���Δf4ȀEf���:`�Gx%X��ʴ�_��L���=��:gYr`!c�������1�� ��� ��ڱL	�=��!���:O
�"�f7T`�/���%axD"�'iw�eH�ŏ%�+���ª��HvKQ5�5�.����}?�Ni=�j�O�۩T$M5Kj�%���[�i����X[�����.i4��a%wn`͉�Sa��q���� [��/�,�4BƇ�`�ԊW���ڍ^�\S�hO��a�X�ʊ)ȇF���8��{���na9�Z�b���|q�~m��>���!@Ր���გ\�1�&L[1vS�<:��(ZBu���4&��ѡ
��'�a"���c��wyu-�����?�%0���K$�R;ߍi�,��r�"0� DGL@yVR�����j��5*������2�\�`��F���(}����Q���ꑄMIϩה�VGm���Y�ʾT2�y�mQR��Љ(dn"�V��.�1���{)s��J1�\L����^v�o���$pp��|�Y�u�L㎇P�3��V��%��W�+?�h�'
�	�R��
�,;,=֘�(� O�e�$��gڕ��%�T
�|%�c�bw�l ed+�n�Cwh��E�s�ka�\���+��G�%ߗJ�J�nKq�),�S�jv��uМJl=�	����a*��e:����Ͳ�(+�5��@��E�����ģڄ����A�os	+е�]��gD��z���9�tP�%�_r���j�\�!`�ԊU&"�`)W�,1%S���1F�6���y��]����&v�$�/���^�m��T���f-�Ё��
{ΚjH-)Zl�A�=��h�@}w��k8<c�4$�_��ag��M?��cG%9Ǥ�;�9�������.#�[��B5d��\�/BvgU�Jl���r&��{��l�}���ux
a~���dB���4Z>��wEV ������j�ܢ�ڮĜԹ�_e�'o���� ��Y�1ڽ�Z�}����~���k8 I9�޺kP:�T���8țZ�ⷍ������ڽ0��<�9�	a��ԝ"ψ7�W����5���Y_Q��D1��N��\�*��GE�,��-I� ��u'������pii-�r��8>��3]�f[�G+�M-�B�k�Օk�I�[�f�j�﯇=<pX�+��9~[��τ$�ȳ����z�M���a��M�7�¿������٬��©ŇzMm8��|]� ���8�j�"@R�&��/&0g ��;�j{d��DJ!��	�@�es������͆�%�р~�W��u�nX�n�י[��ʀp�$K�q~�@��=_V�µW�"e�t����a��>,&�6�!y~�w�3�f�it����b�̀�
sy�	��x&	��v�+����VA��5��o��Z ��7�\e��k��f��� v�|%�7��P�!�vwu;!<X���Ҋ�s���l���qFɏF�6��������9B�<Jڅv��Kп��:q�9�#��7�cΧ�wRZ������f�/��m �h�M��"��� ������C�W�G�C���F@����|��X�'K�
k`�8����v<>��I�c<|ؼ���m��6ZM�c��/����!}"�Vk>(�}
2 *�8$�-��mke��ӣ{�[)�!]en�'�Jq�%Rz�-�O�=0�y0��k��Wynp��}/%�1�A��H��o�K��rk���|/?�(:Eb�Q�\$��L��R(�)j����T~�T%�}́f���j /�b?�14�l�|o)=�ԓ�wK�C5훔���}�MC�F(wB2�Y�zO�]ܬ�VbP�@St9������]����;6͝z�4�~g��#�H�(�9,�G��;��"�ƈAL�a%���� q#�> �K�q*A%�50A�IUQie����_�,:U@�F�~��5��;^��q̡,4fo��A�S����^�v�n�g����vX�ݵ�E���i?�g��ef�:����ṘjgP���!v����o�OC.g!���
�/Y/���Rf?
1z�b`�\Fr���cώ7ߺ�K�743���K�sr������������-��}����Rf/6��ډ� }�<�c�����{�ꤔ�x2�f�J)�$�ٛ�8�ޓ�O��[I�ީ1�g�R��9��^B����&��K@�ܙ�=��I��2r�����q����l���l}t���#��0�Oc�#�wC
>J���:��Q���6�e��K�P�"�h��(Tk�'�s�n2"s �].��a��ȌZ.�tS�f��[�B*�'�u�sY��4ི��J3���3�dߺ*N��"O�_ܪ\��{}�?%H'��rX�7H���i`�9��_�����PU�O�����C�nFYW��ax��j9f�q{���K�����+��f�3���� �*$A�����bِ��t�������<+��"
Lxf4�+Ԭ9�H7{��C������'�H?t-�Hw��g���V���F5���z|��9�@���(j��P|<k�a�N���A�@�=2���!���w�VO[#��'+S0�}$|�Ɛ*_��q�Z��)Sq �{��q���n�Ҳ����Fٽ��1��?ļ*'/��P�J��h_�B�{g9��g��N���(@>)�<�YEb���cAhx�@����ȩ�[�N~_!;��4�jt��K���tDH���=o{Fq���ϻS|���=����1^ӌ��\l��p�r�7�2đ�-@S#S0WQH�ů+`�($��j7��o4�V��s�݄��Wȥ�/������ yb�Xh�{��縰K�Ac֩�&� V9b���%2�iT��Ta����@�L�4Z��B}��fpE�h-̀Y�z����Ы�1I��[e��\��9X F�� ��c�](���|ؒ;�?�-]�K��כ���K}�_��?ۅa���b���C�ك��p�� `��}u�J�0=��:��4��ψ�8����Wү`v*%��E\�w��7
�9�z�ޣ��=L/�5���0�HB�8�0c�F\�~�)���Y�� ;Qƅv�&]a{M���`L~� ����Etl���7R���[������ָ8 F�����S�(Ju]�3��Cj�I�
fR�^�D��%���Ќl��,�NN�)"`Xf�a��`�\��;M����B;:��Q�h�9XܷC:��q�>ˬGN�����Z*o��O�N��Hز���X��M�Lrz	�@\�c�;�S�G}2�O��]uvg��T�p��6J�{�;`�/�:�
A�2Y�R��e���3��vWK�vͧ
@���o�7�C� {�t&M漛�r]g�y�٠e�BF?�w���ܣ���P�V�
f�<�_�Tv���-��r����*�"e�&C���Ӵ�k<��㪦���'K�J�ܹY�/F��^O[rݙі�4����?����wĶ�M�=�����P�}h�p_D�[�4?NE��R~}��� a�;t���y"��%X���V�?�;�o;C��W%�?�H��_��Z��;�o,�P/�wdv�u�W�o��J�����LiƜ����+g��`۝̋��S|!�"Ш($K�/�%T�������/2	z��]�1>&��5�$��+YTY�懻��a���H����:)^B�L��=c�����B"m0)#;k�F�u[E>9Q�kP^���MZ�� �����Y�菺�T_	�
�"��q�b���������ww8�g�t��G��Z�[zؑ���1�nْ?m��&ܽ�IKw�_o�^�7��ߖA�x�1S��GU� 4�&Q1���+�F;E�͡_�0Ao�9��N��AC}�>=+WY�^�F�t�\ke/�}�E���˼���z@5��$+���O�\v�cL����W�^�%i|�F�Xe�z�Sv�K�\D�X���dP��-��ct�� `�t��g8z��fK��d�ͽ�Z(�$��"�=B�#R�i�p��Z�F���T�W������;ԇd��\Z�SL`Y&��[����� ��'���d�k�۫�@�HZ���YxUp���sj!�8��8јꌰX^p�?2h������R�$+(Î�m�1�����K�n�4�����8行�x������:��K/9q<�iiM���v�^��H<^sA��и���cBw�A��?y�Y�M|�s�8��6D�:G�9�CWCn1 [��e��f�'�u65���s���ٮ]���y����[�	��hG�Ǧ��N~K���C_"�/���S������>�Xѕn�u[�ع���2���\�F��^�Op��D��W"�)ӰA���6�r�:2�[��pq�#�f	:Ǥ�1dR�ӂ9�u��8aɋ�P�,�;!�݀l�F*,�����CA+I�Ԝ�団P�I��l�~��NL���"H|DB�c4ʗ�\�sC���B[���������nsʄk�)<�|������>Ęm��sƕ8	��Z�X�PlY
!ɘv��b�-%xb�~��4��O�U' v.b�ԋ��u��l	��͋*ڑ�h��"V��;]zҦ�b��� 4 �ur�
��(ݞ�8۵(e�
�bE��o9�*b�Λ���m6gZ���~Y{pV±����BT��l�Y�0�.�Bek��bb�x�#sws���,r�ʳ �7�cq	��Mi��F�Dcߵb'�ë;)�8]O�ux��O7�Է�����d2��I���@rѢ�|t��?�68�\Ce�]TA�THY0p(f{T�~�9�dl�����̦ &ΎG��P��QC������2�i�9L�`!1�ϓeT�(;�3��zC���M���d����xow/��D���}�[����Đ�n"�v���]��'�veTi�W4U4A�����mnV���F|�Ktk�`�s5A׼�������W<T��v��yF��1x�)���h����Z���mDT P*l���{���XQ����=|P��e�v����r�Qp���6�&7���vdmy�-����YΕ��b�jg8 u��`%�h�7l�cf�u�O1���qu��Ih�F+b����c巀jo����D^dϡ��$��Qo��Lv^�秦�Gɹ�\Uo5XI�1Pȝl�̱��
.Fnmtg'�帥l)�'	g@�
.٫�h����,��PC�n{�<�-�+>�9�L�0��|�ܐ�N�`�;��o�ز�;��;�w�/��Dʛ����z���ok�Gg�]aL�yǼHf��ԧ���2�&I}�0y_�+k�$��p)�Qv���O��:zۿ<�Kg�/g�y���e
��G��D�T>k�q�oG՚�v�I�ݲk|X��f�~�d:V`S�q�M�����K$����K'��:0z7���"�#�7Dy�8_�$(��g؎�
�Y�ə|�_�'8�Įv�YOao�mGg�����m�L� ��@�<1��6T��A��٣t��7"�\�6-[a�y��8�n(�E�`^w��>�Ꮵ���}�����<�B[��-�&��r �*PV8����_}Gr�,:��rp���1삯r�d��x��FI|y��m���}KC�'G|�Oq��b$�>�S}7��:����D��v`���