module testbench_4();

timeunit 10ns;	// Half clock cycle at 50 MHz
			// This is the amount of time represented by #1 
timeprecision 1ns;

// These signals are internal because the processor will be 
// instantiated as a submodule in testbench.
logic Clk = 0;
logic Reset, ClearA_LoadB, Run;
logic [7:0] S;
logic 		X;
logic [7:0] Aval,Bval;
logic [6:0] AhexL,
		 AhexU,
		 BhexL,
		 BhexU; 

				
// A counter to count the instances where simulation results
// do no match with expected results
//integer ErrorCnt = 0;
		
// Instantiating the DUT
// Make sure the module and signal names match with those in your design
lab4_8_bit_multiplier_toplevel mt(.*);

// Toggle the clock
// #1 means wait for a delay of 1 timeunit
always begin : CLOCK_GENERATION
#1 Clk = ~Clk;
end

initial begin: CLOCK_INITIALIZATION
    Clk = 0;
end 

// Testing begins here
// The initial block is not synthesizable
// Everything happens sequentially inside an initial block
// as in a software program
initial begin: TEST_VECTORS
Reset = 0;		// Toggle loadB clearA
ClearA_LoadB = 1;
Run = 1;
S = 8'b00000011;
//S = 8'h1;	// Specify S --load into B


#2 ClearA_LoadB = 0;
Reset = 1;

#4 ClearA_LoadB = 1;
	Run = 0;	
#22;
end

endmodule
